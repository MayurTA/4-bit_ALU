magic
tech scmos
timestamp 1607684136
<< ab >>
rect 3 232 4 240
rect 6 168 30 240
rect 32 232 63 240
rect 39 193 63 232
rect 78 205 134 240
rect 136 232 143 240
rect 78 201 132 205
rect 39 189 67 193
rect 32 168 37 176
rect 39 168 63 189
rect 78 176 134 201
rect 144 193 166 240
rect 142 189 166 193
rect 144 176 166 189
rect 65 168 134 176
rect 136 168 143 176
rect 144 168 175 176
rect 176 168 200 240
rect 202 232 208 240
rect 210 232 313 240
rect 314 232 384 240
rect 210 168 274 232
rect 281 176 313 232
rect 276 169 313 176
rect 320 173 384 232
rect 320 169 386 173
rect 276 168 353 169
rect 355 168 386 169
rect 388 168 428 240
rect 430 232 438 240
rect 440 168 480 240
rect 482 168 522 240
rect 526 168 566 240
rect 5 115 230 168
rect 231 160 244 168
rect 245 115 470 168
rect 471 160 479 168
rect 482 167 485 168
rect 5 110 233 115
rect 245 110 473 115
rect 5 82 230 110
rect 245 104 470 110
rect 502 104 566 168
rect 231 97 470 104
rect 471 97 479 104
rect 480 97 566 104
rect 231 96 566 97
rect 231 88 242 96
rect 244 82 469 96
rect 2 77 230 82
rect 241 77 469 82
rect 4 58 230 77
rect 5 -29 230 58
rect 231 24 242 32
rect 244 24 469 77
rect 470 88 566 96
rect 470 64 485 88
rect 502 64 566 88
rect 503 32 566 64
rect 470 24 566 32
rect 231 16 244 24
rect 245 23 500 24
rect 245 -29 470 23
rect 471 16 479 23
rect 485 16 500 23
rect 5 -34 233 -29
rect 245 -34 473 -29
rect 5 -62 230 -34
rect 245 -40 470 -34
rect 231 -47 470 -40
rect 471 -47 479 -40
rect 480 -47 485 -40
rect 231 -48 485 -47
rect 231 -56 242 -48
rect 244 -62 469 -48
rect 2 -67 230 -62
rect 241 -67 469 -62
rect 5 -120 230 -67
rect 231 -120 242 -112
rect 244 -120 469 -67
rect 470 -80 485 -48
rect 470 -120 501 -112
rect 502 -120 566 24
<< nwell >>
rect 0 128 571 208
rect 0 -16 571 64
rect 0 -125 571 -80
<< pwell >>
rect 0 208 571 245
rect 0 64 571 128
rect 0 -80 571 -16
<< poly >>
rect 19 228 21 233
rect 52 228 54 233
rect 93 227 95 232
rect 103 227 105 232
rect 219 236 238 238
rect 113 225 115 229
rect 123 225 125 229
rect 153 228 155 233
rect 189 228 191 233
rect 219 228 221 236
rect 229 228 231 232
rect 236 228 238 236
rect 329 236 348 238
rect 246 228 248 233
rect 253 228 255 233
rect 263 228 265 233
rect 302 231 304 236
rect 19 211 21 214
rect 52 211 54 214
rect 14 209 21 211
rect 14 207 16 209
rect 18 207 21 209
rect 14 205 21 207
rect 47 209 54 211
rect 47 207 49 209
rect 51 207 54 209
rect 47 205 54 207
rect 93 205 95 221
rect 103 218 105 221
rect 99 216 105 218
rect 99 214 101 216
rect 103 214 105 216
rect 99 212 105 214
rect 19 202 21 205
rect 52 202 54 205
rect 87 203 95 205
rect 87 201 89 203
rect 91 201 95 203
rect 87 199 95 201
rect 93 196 95 199
rect 100 196 102 212
rect 113 211 115 219
rect 109 209 115 211
rect 109 208 111 209
rect 107 207 111 208
rect 113 207 115 209
rect 107 205 115 207
rect 123 205 125 219
rect 292 225 294 230
rect 107 196 109 205
rect 119 203 125 205
rect 119 201 121 203
rect 123 201 125 203
rect 153 211 155 214
rect 189 211 191 214
rect 153 209 160 211
rect 153 207 156 209
rect 158 207 160 209
rect 153 205 160 207
rect 184 209 191 211
rect 184 207 186 209
rect 188 207 191 209
rect 184 205 191 207
rect 153 202 155 205
rect 189 202 191 205
rect 219 202 221 222
rect 229 211 231 222
rect 225 209 231 211
rect 225 207 227 209
rect 229 207 231 209
rect 236 209 238 222
rect 246 219 248 222
rect 242 217 248 219
rect 242 215 244 217
rect 246 215 248 217
rect 242 213 248 215
rect 253 209 255 222
rect 263 219 265 222
rect 260 217 266 219
rect 260 215 262 217
rect 264 215 266 217
rect 260 213 266 215
rect 329 228 331 236
rect 339 228 341 232
rect 346 228 348 236
rect 356 228 358 233
rect 363 228 365 233
rect 373 228 375 233
rect 397 229 399 234
rect 407 229 409 234
rect 417 229 419 234
rect 449 229 451 234
rect 459 229 461 234
rect 469 229 471 234
rect 491 229 493 234
rect 501 229 503 234
rect 511 229 513 234
rect 535 229 537 234
rect 545 229 547 234
rect 555 229 557 234
rect 236 207 248 209
rect 225 205 231 207
rect 114 199 125 201
rect 114 196 116 199
rect 19 170 21 174
rect 52 170 54 174
rect 93 170 95 174
rect 100 170 102 174
rect 107 170 109 174
rect 114 170 116 174
rect 219 193 221 196
rect 212 191 221 193
rect 229 194 231 205
rect 235 201 241 203
rect 235 199 237 201
rect 239 199 241 201
rect 235 197 241 199
rect 236 194 238 197
rect 246 194 248 207
rect 252 207 258 209
rect 252 205 254 207
rect 256 205 258 207
rect 252 203 258 205
rect 253 194 255 203
rect 263 194 265 213
rect 292 211 294 214
rect 302 211 304 214
rect 291 209 304 211
rect 291 207 293 209
rect 295 207 304 209
rect 291 205 304 207
rect 292 202 294 205
rect 302 202 304 205
rect 329 202 331 222
rect 339 211 341 222
rect 335 209 341 211
rect 335 207 337 209
rect 339 207 341 209
rect 346 209 348 222
rect 356 219 358 222
rect 352 217 358 219
rect 352 215 354 217
rect 356 215 358 217
rect 352 213 358 215
rect 363 209 365 222
rect 373 219 375 222
rect 370 217 376 219
rect 370 215 372 217
rect 374 215 376 217
rect 370 213 376 215
rect 346 207 358 209
rect 335 205 341 207
rect 212 189 214 191
rect 216 189 218 191
rect 212 187 218 189
rect 229 177 231 182
rect 236 177 238 182
rect 246 177 248 182
rect 253 177 255 182
rect 263 177 265 182
rect 153 170 155 174
rect 189 170 191 174
rect 329 193 331 196
rect 322 191 331 193
rect 339 194 341 205
rect 345 201 351 203
rect 345 199 347 201
rect 349 199 351 201
rect 345 197 351 199
rect 346 194 348 197
rect 356 194 358 207
rect 362 207 368 209
rect 362 205 364 207
rect 366 205 368 207
rect 362 203 368 205
rect 363 194 365 203
rect 373 194 375 213
rect 397 211 399 215
rect 407 212 409 215
rect 417 212 419 215
rect 396 209 402 211
rect 396 207 398 209
rect 400 207 402 209
rect 396 205 402 207
rect 406 210 419 212
rect 449 211 451 215
rect 459 212 461 215
rect 469 212 471 215
rect 406 208 408 210
rect 410 208 419 210
rect 406 206 419 208
rect 397 202 399 205
rect 407 202 409 206
rect 417 202 419 206
rect 448 209 454 211
rect 448 207 450 209
rect 452 207 454 209
rect 448 205 454 207
rect 458 210 471 212
rect 491 211 493 215
rect 501 212 503 215
rect 511 212 513 215
rect 458 208 460 210
rect 462 208 471 210
rect 458 206 471 208
rect 449 202 451 205
rect 459 202 461 206
rect 469 202 471 206
rect 490 209 496 211
rect 490 207 492 209
rect 494 207 496 209
rect 490 205 496 207
rect 500 210 513 212
rect 535 211 537 215
rect 545 212 547 215
rect 555 212 557 215
rect 500 208 502 210
rect 504 208 513 210
rect 500 206 513 208
rect 491 202 493 205
rect 501 202 503 206
rect 511 202 513 206
rect 534 209 540 211
rect 534 207 536 209
rect 538 207 540 209
rect 534 205 540 207
rect 544 210 557 212
rect 544 208 546 210
rect 548 208 557 210
rect 544 206 557 208
rect 535 202 537 205
rect 545 202 547 206
rect 555 202 557 206
rect 322 189 324 191
rect 326 189 328 191
rect 322 187 328 189
rect 339 177 341 182
rect 346 177 348 182
rect 356 177 358 182
rect 363 177 365 182
rect 373 177 375 182
rect 292 170 294 174
rect 302 170 304 174
rect 397 170 399 174
rect 407 170 409 174
rect 417 170 419 174
rect 449 170 451 174
rect 459 170 461 174
rect 469 170 471 174
rect 491 170 493 174
rect 501 170 503 174
rect 511 170 513 174
rect 535 170 537 174
rect 545 170 547 174
rect 555 170 557 174
rect 14 162 16 166
rect 37 159 39 164
rect 44 159 46 164
rect 62 162 64 166
rect 72 162 74 166
rect 82 162 84 166
rect 110 162 112 166
rect 27 150 29 155
rect 14 124 16 137
rect 27 134 29 137
rect 133 159 135 164
rect 140 159 142 164
rect 158 162 160 166
rect 168 162 170 166
rect 178 162 180 166
rect 199 162 201 166
rect 206 162 208 166
rect 123 150 125 155
rect 20 132 29 134
rect 20 130 22 132
rect 24 130 26 132
rect 37 131 39 134
rect 44 131 46 134
rect 62 131 64 134
rect 72 131 74 134
rect 82 131 84 134
rect 20 128 26 130
rect 14 122 20 124
rect 14 120 16 122
rect 18 120 20 122
rect 14 118 20 120
rect 14 115 16 118
rect 24 115 26 128
rect 34 129 40 131
rect 34 127 36 129
rect 38 127 40 129
rect 34 125 40 127
rect 44 129 66 131
rect 44 127 55 129
rect 57 127 62 129
rect 64 127 66 129
rect 44 125 66 127
rect 70 129 76 131
rect 70 127 72 129
rect 74 127 76 129
rect 70 125 76 127
rect 80 129 86 131
rect 80 127 82 129
rect 84 127 86 129
rect 80 125 86 127
rect 34 122 36 125
rect 44 122 46 125
rect 64 122 66 125
rect 71 122 73 125
rect 14 98 16 102
rect 24 100 26 105
rect 34 103 36 108
rect 44 103 46 108
rect 82 116 84 125
rect 110 124 112 137
rect 123 134 125 137
rect 219 162 221 166
rect 254 162 256 166
rect 277 159 279 164
rect 284 159 286 164
rect 302 162 304 166
rect 312 162 314 166
rect 322 162 324 166
rect 350 162 352 166
rect 267 150 269 155
rect 116 132 125 134
rect 116 130 118 132
rect 120 130 122 132
rect 133 131 135 134
rect 140 131 142 134
rect 158 131 160 134
rect 168 131 170 134
rect 178 131 180 134
rect 199 131 201 134
rect 206 131 208 134
rect 219 131 221 134
rect 116 128 122 130
rect 110 122 116 124
rect 110 120 112 122
rect 114 120 116 122
rect 110 118 116 120
rect 110 115 112 118
rect 120 115 122 128
rect 130 129 136 131
rect 130 127 132 129
rect 134 127 136 129
rect 130 125 136 127
rect 140 129 162 131
rect 140 127 151 129
rect 153 127 158 129
rect 160 127 162 129
rect 140 125 162 127
rect 166 129 172 131
rect 166 127 168 129
rect 170 127 172 129
rect 166 125 172 127
rect 176 129 182 131
rect 176 127 178 129
rect 180 127 182 129
rect 176 125 182 127
rect 192 129 201 131
rect 192 127 194 129
rect 196 127 201 129
rect 192 125 201 127
rect 205 129 211 131
rect 205 127 207 129
rect 209 127 211 129
rect 205 125 211 127
rect 215 129 221 131
rect 215 127 217 129
rect 219 127 221 129
rect 215 125 221 127
rect 130 122 132 125
rect 140 122 142 125
rect 160 122 162 125
rect 167 122 169 125
rect 64 98 66 102
rect 71 98 73 102
rect 82 98 84 102
rect 110 98 112 102
rect 120 100 122 105
rect 130 103 132 108
rect 140 103 142 108
rect 178 116 180 125
rect 199 119 201 125
rect 209 117 211 125
rect 219 122 221 125
rect 254 124 256 137
rect 267 134 269 137
rect 373 159 375 164
rect 380 159 382 164
rect 398 162 400 166
rect 408 162 410 166
rect 418 162 420 166
rect 439 162 441 166
rect 446 162 448 166
rect 363 150 365 155
rect 260 132 269 134
rect 260 130 262 132
rect 264 130 266 132
rect 277 131 279 134
rect 284 131 286 134
rect 302 131 304 134
rect 312 131 314 134
rect 322 131 324 134
rect 260 128 266 130
rect 254 122 260 124
rect 199 107 201 111
rect 209 104 211 109
rect 254 120 256 122
rect 258 120 260 122
rect 254 118 260 120
rect 254 115 256 118
rect 264 115 266 128
rect 274 129 280 131
rect 274 127 276 129
rect 278 127 280 129
rect 274 125 280 127
rect 284 129 306 131
rect 284 127 295 129
rect 297 127 302 129
rect 304 127 306 129
rect 284 125 306 127
rect 310 129 316 131
rect 310 127 312 129
rect 314 127 316 129
rect 310 125 316 127
rect 320 129 326 131
rect 320 127 322 129
rect 324 127 326 129
rect 320 125 326 127
rect 274 122 276 125
rect 284 122 286 125
rect 304 122 306 125
rect 311 122 313 125
rect 219 103 221 108
rect 160 98 162 102
rect 167 98 169 102
rect 178 98 180 102
rect 254 98 256 102
rect 264 100 266 105
rect 274 103 276 108
rect 284 103 286 108
rect 322 116 324 125
rect 350 124 352 137
rect 363 134 365 137
rect 459 162 461 166
rect 521 154 523 159
rect 528 154 530 159
rect 538 154 540 159
rect 545 154 547 159
rect 555 154 557 159
rect 504 147 510 149
rect 504 145 506 147
rect 508 145 510 147
rect 504 143 513 145
rect 511 140 513 143
rect 356 132 365 134
rect 356 130 358 132
rect 360 130 362 132
rect 373 131 375 134
rect 380 131 382 134
rect 398 131 400 134
rect 408 131 410 134
rect 418 131 420 134
rect 439 131 441 134
rect 446 131 448 134
rect 459 131 461 134
rect 356 128 362 130
rect 350 122 356 124
rect 350 120 352 122
rect 354 120 356 122
rect 350 118 356 120
rect 350 115 352 118
rect 360 115 362 128
rect 370 129 376 131
rect 370 127 372 129
rect 374 127 376 129
rect 370 125 376 127
rect 380 129 402 131
rect 380 127 391 129
rect 393 127 398 129
rect 400 127 402 129
rect 380 125 402 127
rect 406 129 412 131
rect 406 127 408 129
rect 410 127 412 129
rect 406 125 412 127
rect 416 129 422 131
rect 416 127 418 129
rect 420 127 422 129
rect 416 125 422 127
rect 432 129 441 131
rect 432 127 434 129
rect 436 127 441 129
rect 432 125 441 127
rect 445 129 451 131
rect 445 127 447 129
rect 449 127 451 129
rect 445 125 451 127
rect 455 129 461 131
rect 455 127 457 129
rect 459 127 461 129
rect 455 125 461 127
rect 370 122 372 125
rect 380 122 382 125
rect 400 122 402 125
rect 407 122 409 125
rect 304 98 306 102
rect 311 98 313 102
rect 322 98 324 102
rect 350 98 352 102
rect 360 100 362 105
rect 370 103 372 108
rect 380 103 382 108
rect 418 116 420 125
rect 439 119 441 125
rect 449 117 451 125
rect 459 122 461 125
rect 439 107 441 111
rect 449 104 451 109
rect 511 114 513 134
rect 521 131 523 142
rect 528 139 530 142
rect 527 137 533 139
rect 527 135 529 137
rect 531 135 533 137
rect 527 133 533 135
rect 517 129 523 131
rect 538 129 540 142
rect 545 133 547 142
rect 517 127 519 129
rect 521 127 523 129
rect 517 125 523 127
rect 521 114 523 125
rect 528 127 540 129
rect 544 131 550 133
rect 544 129 546 131
rect 548 129 550 131
rect 544 127 550 129
rect 528 114 530 127
rect 534 121 540 123
rect 534 119 536 121
rect 538 119 540 121
rect 534 117 540 119
rect 538 114 540 117
rect 545 114 547 127
rect 555 123 557 142
rect 552 121 558 123
rect 552 119 554 121
rect 556 119 558 121
rect 552 117 558 119
rect 555 114 557 117
rect 459 103 461 108
rect 400 98 402 102
rect 407 98 409 102
rect 418 98 420 102
rect 511 100 513 108
rect 521 104 523 108
rect 528 100 530 108
rect 538 103 540 108
rect 545 103 547 108
rect 555 103 557 108
rect 511 98 530 100
rect 55 90 57 94
rect 66 90 68 94
rect 73 90 75 94
rect 14 84 16 89
rect 24 83 26 88
rect 34 81 36 85
rect 14 67 16 70
rect 24 67 26 75
rect 34 67 36 73
rect 55 67 57 76
rect 93 84 95 89
rect 103 84 105 89
rect 113 87 115 92
rect 123 90 125 94
rect 151 90 153 94
rect 162 90 164 94
rect 169 90 171 94
rect 66 67 68 70
rect 73 67 75 70
rect 93 67 95 70
rect 103 67 105 70
rect 14 65 20 67
rect 14 63 16 65
rect 18 63 20 65
rect 14 61 20 63
rect 24 65 30 67
rect 24 63 26 65
rect 28 63 30 65
rect 24 61 30 63
rect 34 65 43 67
rect 34 63 39 65
rect 41 63 43 65
rect 34 61 43 63
rect 53 65 59 67
rect 53 63 55 65
rect 57 63 59 65
rect 53 61 59 63
rect 63 65 69 67
rect 63 63 65 65
rect 67 63 69 65
rect 63 61 69 63
rect 73 65 95 67
rect 73 63 75 65
rect 77 63 82 65
rect 84 63 95 65
rect 73 61 95 63
rect 99 65 105 67
rect 99 63 101 65
rect 103 63 105 65
rect 99 61 105 63
rect 113 64 115 77
rect 123 74 125 77
rect 119 72 125 74
rect 119 70 121 72
rect 123 70 125 72
rect 119 68 125 70
rect 113 62 119 64
rect 14 58 16 61
rect 27 58 29 61
rect 34 58 36 61
rect 55 58 57 61
rect 65 58 67 61
rect 75 58 77 61
rect 93 58 95 61
rect 100 58 102 61
rect 113 60 115 62
rect 117 60 119 62
rect 110 58 119 60
rect 14 26 16 30
rect 110 55 112 58
rect 123 55 125 68
rect 151 67 153 76
rect 189 84 191 89
rect 199 84 201 89
rect 209 87 211 92
rect 219 90 221 94
rect 294 90 296 94
rect 305 90 307 94
rect 312 90 314 94
rect 253 84 255 89
rect 162 67 164 70
rect 169 67 171 70
rect 189 67 191 70
rect 199 67 201 70
rect 149 65 155 67
rect 149 63 151 65
rect 153 63 155 65
rect 149 61 155 63
rect 159 65 165 67
rect 159 63 161 65
rect 163 63 165 65
rect 159 61 165 63
rect 169 65 191 67
rect 169 63 171 65
rect 173 63 178 65
rect 180 63 191 65
rect 169 61 191 63
rect 195 65 201 67
rect 195 63 197 65
rect 199 63 201 65
rect 195 61 201 63
rect 209 64 211 77
rect 219 74 221 77
rect 215 72 221 74
rect 215 70 217 72
rect 219 70 221 72
rect 263 83 265 88
rect 273 81 275 85
rect 215 68 221 70
rect 209 62 215 64
rect 151 58 153 61
rect 161 58 163 61
rect 171 58 173 61
rect 189 58 191 61
rect 196 58 198 61
rect 209 60 211 62
rect 213 60 215 62
rect 206 58 215 60
rect 110 37 112 42
rect 27 26 29 30
rect 34 26 36 30
rect 55 26 57 30
rect 65 26 67 30
rect 75 26 77 30
rect 93 28 95 33
rect 100 28 102 33
rect 206 55 208 58
rect 219 55 221 68
rect 253 67 255 70
rect 263 67 265 75
rect 273 67 275 73
rect 294 67 296 76
rect 332 84 334 89
rect 342 84 344 89
rect 352 87 354 92
rect 362 90 364 94
rect 390 90 392 94
rect 401 90 403 94
rect 408 90 410 94
rect 305 67 307 70
rect 312 67 314 70
rect 332 67 334 70
rect 342 67 344 70
rect 253 65 259 67
rect 253 63 255 65
rect 257 63 259 65
rect 253 61 259 63
rect 263 65 269 67
rect 263 63 265 65
rect 267 63 269 65
rect 263 61 269 63
rect 273 65 282 67
rect 273 63 278 65
rect 280 63 282 65
rect 273 61 282 63
rect 292 65 298 67
rect 292 63 294 65
rect 296 63 298 65
rect 292 61 298 63
rect 302 65 308 67
rect 302 63 304 65
rect 306 63 308 65
rect 302 61 308 63
rect 312 65 334 67
rect 312 63 314 65
rect 316 63 321 65
rect 323 63 334 65
rect 312 61 334 63
rect 338 65 344 67
rect 338 63 340 65
rect 342 63 344 65
rect 338 61 344 63
rect 352 64 354 77
rect 362 74 364 77
rect 358 72 364 74
rect 358 70 360 72
rect 362 70 364 72
rect 358 68 364 70
rect 352 62 358 64
rect 253 58 255 61
rect 266 58 268 61
rect 273 58 275 61
rect 294 58 296 61
rect 304 58 306 61
rect 314 58 316 61
rect 332 58 334 61
rect 339 58 341 61
rect 352 60 354 62
rect 356 60 358 62
rect 349 58 358 60
rect 206 37 208 42
rect 123 26 125 30
rect 151 26 153 30
rect 161 26 163 30
rect 171 26 173 30
rect 189 28 191 33
rect 196 28 198 33
rect 219 26 221 30
rect 253 26 255 30
rect 349 55 351 58
rect 362 55 364 68
rect 390 67 392 76
rect 428 84 430 89
rect 438 84 440 89
rect 448 87 450 92
rect 458 90 460 94
rect 511 92 530 94
rect 511 84 513 92
rect 521 84 523 88
rect 528 84 530 92
rect 538 84 540 89
rect 545 84 547 89
rect 555 84 557 89
rect 401 67 403 70
rect 408 67 410 70
rect 428 67 430 70
rect 438 67 440 70
rect 388 65 394 67
rect 388 63 390 65
rect 392 63 394 65
rect 388 61 394 63
rect 398 65 404 67
rect 398 63 400 65
rect 402 63 404 65
rect 398 61 404 63
rect 408 65 430 67
rect 408 63 410 65
rect 412 63 417 65
rect 419 63 430 65
rect 408 61 430 63
rect 434 65 440 67
rect 434 63 436 65
rect 438 63 440 65
rect 434 61 440 63
rect 448 64 450 77
rect 458 74 460 77
rect 454 72 460 74
rect 454 70 456 72
rect 458 70 460 72
rect 454 68 460 70
rect 448 62 454 64
rect 390 58 392 61
rect 400 58 402 61
rect 410 58 412 61
rect 428 58 430 61
rect 435 58 437 61
rect 448 60 450 62
rect 452 60 454 62
rect 445 58 454 60
rect 349 37 351 42
rect 266 26 268 30
rect 273 26 275 30
rect 294 26 296 30
rect 304 26 306 30
rect 314 26 316 30
rect 332 28 334 33
rect 339 28 341 33
rect 445 55 447 58
rect 458 55 460 68
rect 511 58 513 78
rect 521 67 523 78
rect 517 65 523 67
rect 517 63 519 65
rect 521 63 523 65
rect 528 65 530 78
rect 538 75 540 78
rect 534 73 540 75
rect 534 71 536 73
rect 538 71 540 73
rect 534 69 540 71
rect 545 65 547 78
rect 555 75 557 78
rect 552 73 558 75
rect 552 71 554 73
rect 556 71 558 73
rect 552 69 558 71
rect 528 63 540 65
rect 517 61 523 63
rect 445 37 447 42
rect 362 26 364 30
rect 390 26 392 30
rect 400 26 402 30
rect 410 26 412 30
rect 428 28 430 33
rect 435 28 437 33
rect 511 49 513 52
rect 504 47 513 49
rect 521 50 523 61
rect 527 57 533 59
rect 527 55 529 57
rect 531 55 533 57
rect 527 53 533 55
rect 528 50 530 53
rect 538 50 540 63
rect 544 63 550 65
rect 544 61 546 63
rect 548 61 550 63
rect 544 59 550 61
rect 545 50 547 59
rect 555 50 557 69
rect 504 45 506 47
rect 508 45 510 47
rect 504 43 510 45
rect 521 33 523 38
rect 528 33 530 38
rect 538 33 540 38
rect 545 33 547 38
rect 555 33 557 38
rect 458 26 460 30
rect 14 18 16 22
rect 37 15 39 20
rect 44 15 46 20
rect 62 18 64 22
rect 72 18 74 22
rect 82 18 84 22
rect 110 18 112 22
rect 27 6 29 11
rect 14 -20 16 -7
rect 27 -10 29 -7
rect 133 15 135 20
rect 140 15 142 20
rect 158 18 160 22
rect 168 18 170 22
rect 178 18 180 22
rect 199 18 201 22
rect 206 18 208 22
rect 123 6 125 11
rect 20 -12 29 -10
rect 20 -14 22 -12
rect 24 -14 26 -12
rect 37 -13 39 -10
rect 44 -13 46 -10
rect 62 -13 64 -10
rect 72 -13 74 -10
rect 82 -13 84 -10
rect 20 -16 26 -14
rect 14 -22 20 -20
rect 14 -24 16 -22
rect 18 -24 20 -22
rect 14 -26 20 -24
rect 14 -29 16 -26
rect 24 -29 26 -16
rect 34 -15 40 -13
rect 34 -17 36 -15
rect 38 -17 40 -15
rect 34 -19 40 -17
rect 44 -15 66 -13
rect 44 -17 55 -15
rect 57 -17 62 -15
rect 64 -17 66 -15
rect 44 -19 66 -17
rect 70 -15 76 -13
rect 70 -17 72 -15
rect 74 -17 76 -15
rect 70 -19 76 -17
rect 80 -15 86 -13
rect 80 -17 82 -15
rect 84 -17 86 -15
rect 80 -19 86 -17
rect 34 -22 36 -19
rect 44 -22 46 -19
rect 64 -22 66 -19
rect 71 -22 73 -19
rect 14 -46 16 -42
rect 24 -44 26 -39
rect 34 -41 36 -36
rect 44 -41 46 -36
rect 82 -28 84 -19
rect 110 -20 112 -7
rect 123 -10 125 -7
rect 219 18 221 22
rect 254 18 256 22
rect 277 15 279 20
rect 284 15 286 20
rect 302 18 304 22
rect 312 18 314 22
rect 322 18 324 22
rect 350 18 352 22
rect 267 6 269 11
rect 116 -12 125 -10
rect 116 -14 118 -12
rect 120 -14 122 -12
rect 133 -13 135 -10
rect 140 -13 142 -10
rect 158 -13 160 -10
rect 168 -13 170 -10
rect 178 -13 180 -10
rect 199 -13 201 -10
rect 206 -13 208 -10
rect 219 -13 221 -10
rect 116 -16 122 -14
rect 110 -22 116 -20
rect 110 -24 112 -22
rect 114 -24 116 -22
rect 110 -26 116 -24
rect 110 -29 112 -26
rect 120 -29 122 -16
rect 130 -15 136 -13
rect 130 -17 132 -15
rect 134 -17 136 -15
rect 130 -19 136 -17
rect 140 -15 162 -13
rect 140 -17 151 -15
rect 153 -17 158 -15
rect 160 -17 162 -15
rect 140 -19 162 -17
rect 166 -15 172 -13
rect 166 -17 168 -15
rect 170 -17 172 -15
rect 166 -19 172 -17
rect 176 -15 182 -13
rect 176 -17 178 -15
rect 180 -17 182 -15
rect 176 -19 182 -17
rect 192 -15 201 -13
rect 192 -17 194 -15
rect 196 -17 201 -15
rect 192 -19 201 -17
rect 205 -15 211 -13
rect 205 -17 207 -15
rect 209 -17 211 -15
rect 205 -19 211 -17
rect 215 -15 221 -13
rect 215 -17 217 -15
rect 219 -17 221 -15
rect 215 -19 221 -17
rect 130 -22 132 -19
rect 140 -22 142 -19
rect 160 -22 162 -19
rect 167 -22 169 -19
rect 64 -46 66 -42
rect 71 -46 73 -42
rect 82 -46 84 -42
rect 110 -46 112 -42
rect 120 -44 122 -39
rect 130 -41 132 -36
rect 140 -41 142 -36
rect 178 -28 180 -19
rect 199 -25 201 -19
rect 209 -27 211 -19
rect 219 -22 221 -19
rect 254 -20 256 -7
rect 267 -10 269 -7
rect 373 15 375 20
rect 380 15 382 20
rect 398 18 400 22
rect 408 18 410 22
rect 418 18 420 22
rect 439 18 441 22
rect 446 18 448 22
rect 363 6 365 11
rect 260 -12 269 -10
rect 260 -14 262 -12
rect 264 -14 266 -12
rect 277 -13 279 -10
rect 284 -13 286 -10
rect 302 -13 304 -10
rect 312 -13 314 -10
rect 322 -13 324 -10
rect 260 -16 266 -14
rect 254 -22 260 -20
rect 199 -37 201 -33
rect 209 -40 211 -35
rect 254 -24 256 -22
rect 258 -24 260 -22
rect 254 -26 260 -24
rect 254 -29 256 -26
rect 264 -29 266 -16
rect 274 -15 280 -13
rect 274 -17 276 -15
rect 278 -17 280 -15
rect 274 -19 280 -17
rect 284 -15 306 -13
rect 284 -17 295 -15
rect 297 -17 302 -15
rect 304 -17 306 -15
rect 284 -19 306 -17
rect 310 -15 316 -13
rect 310 -17 312 -15
rect 314 -17 316 -15
rect 310 -19 316 -17
rect 320 -15 326 -13
rect 320 -17 322 -15
rect 324 -17 326 -15
rect 320 -19 326 -17
rect 274 -22 276 -19
rect 284 -22 286 -19
rect 304 -22 306 -19
rect 311 -22 313 -19
rect 219 -41 221 -36
rect 160 -46 162 -42
rect 167 -46 169 -42
rect 178 -46 180 -42
rect 254 -46 256 -42
rect 264 -44 266 -39
rect 274 -41 276 -36
rect 284 -41 286 -36
rect 322 -28 324 -19
rect 350 -20 352 -7
rect 363 -10 365 -7
rect 459 18 461 22
rect 521 10 523 15
rect 528 10 530 15
rect 538 10 540 15
rect 545 10 547 15
rect 555 10 557 15
rect 504 3 510 5
rect 504 1 506 3
rect 508 1 510 3
rect 504 -1 513 1
rect 511 -4 513 -1
rect 356 -12 365 -10
rect 356 -14 358 -12
rect 360 -14 362 -12
rect 373 -13 375 -10
rect 380 -13 382 -10
rect 398 -13 400 -10
rect 408 -13 410 -10
rect 418 -13 420 -10
rect 439 -13 441 -10
rect 446 -13 448 -10
rect 459 -13 461 -10
rect 356 -16 362 -14
rect 350 -22 356 -20
rect 350 -24 352 -22
rect 354 -24 356 -22
rect 350 -26 356 -24
rect 350 -29 352 -26
rect 360 -29 362 -16
rect 370 -15 376 -13
rect 370 -17 372 -15
rect 374 -17 376 -15
rect 370 -19 376 -17
rect 380 -15 402 -13
rect 380 -17 391 -15
rect 393 -17 398 -15
rect 400 -17 402 -15
rect 380 -19 402 -17
rect 406 -15 412 -13
rect 406 -17 408 -15
rect 410 -17 412 -15
rect 406 -19 412 -17
rect 416 -15 422 -13
rect 416 -17 418 -15
rect 420 -17 422 -15
rect 416 -19 422 -17
rect 432 -15 441 -13
rect 432 -17 434 -15
rect 436 -17 441 -15
rect 432 -19 441 -17
rect 445 -15 451 -13
rect 445 -17 447 -15
rect 449 -17 451 -15
rect 445 -19 451 -17
rect 455 -15 461 -13
rect 455 -17 457 -15
rect 459 -17 461 -15
rect 455 -19 461 -17
rect 370 -22 372 -19
rect 380 -22 382 -19
rect 400 -22 402 -19
rect 407 -22 409 -19
rect 304 -46 306 -42
rect 311 -46 313 -42
rect 322 -46 324 -42
rect 350 -46 352 -42
rect 360 -44 362 -39
rect 370 -41 372 -36
rect 380 -41 382 -36
rect 418 -28 420 -19
rect 439 -25 441 -19
rect 449 -27 451 -19
rect 459 -22 461 -19
rect 439 -37 441 -33
rect 449 -40 451 -35
rect 511 -30 513 -10
rect 521 -13 523 -2
rect 528 -5 530 -2
rect 527 -7 533 -5
rect 527 -9 529 -7
rect 531 -9 533 -7
rect 527 -11 533 -9
rect 517 -15 523 -13
rect 538 -15 540 -2
rect 545 -11 547 -2
rect 517 -17 519 -15
rect 521 -17 523 -15
rect 517 -19 523 -17
rect 521 -30 523 -19
rect 528 -17 540 -15
rect 544 -13 550 -11
rect 544 -15 546 -13
rect 548 -15 550 -13
rect 544 -17 550 -15
rect 528 -30 530 -17
rect 534 -23 540 -21
rect 534 -25 536 -23
rect 538 -25 540 -23
rect 534 -27 540 -25
rect 538 -30 540 -27
rect 545 -30 547 -17
rect 555 -21 557 -2
rect 552 -23 558 -21
rect 552 -25 554 -23
rect 556 -25 558 -23
rect 552 -27 558 -25
rect 555 -30 557 -27
rect 459 -41 461 -36
rect 400 -46 402 -42
rect 407 -46 409 -42
rect 418 -46 420 -42
rect 511 -44 513 -36
rect 521 -40 523 -36
rect 528 -44 530 -36
rect 538 -41 540 -36
rect 545 -41 547 -36
rect 555 -41 557 -36
rect 511 -46 530 -44
rect 55 -54 57 -50
rect 66 -54 68 -50
rect 73 -54 75 -50
rect 14 -60 16 -55
rect 24 -61 26 -56
rect 34 -63 36 -59
rect 14 -77 16 -74
rect 24 -77 26 -69
rect 34 -77 36 -71
rect 55 -77 57 -68
rect 93 -60 95 -55
rect 103 -60 105 -55
rect 113 -57 115 -52
rect 123 -54 125 -50
rect 151 -54 153 -50
rect 162 -54 164 -50
rect 169 -54 171 -50
rect 66 -77 68 -74
rect 73 -77 75 -74
rect 93 -77 95 -74
rect 103 -77 105 -74
rect 14 -79 20 -77
rect 14 -81 16 -79
rect 18 -81 20 -79
rect 14 -83 20 -81
rect 24 -79 30 -77
rect 24 -81 26 -79
rect 28 -81 30 -79
rect 24 -83 30 -81
rect 34 -79 43 -77
rect 34 -81 39 -79
rect 41 -81 43 -79
rect 34 -83 43 -81
rect 53 -79 59 -77
rect 53 -81 55 -79
rect 57 -81 59 -79
rect 53 -83 59 -81
rect 63 -79 69 -77
rect 63 -81 65 -79
rect 67 -81 69 -79
rect 63 -83 69 -81
rect 73 -79 95 -77
rect 73 -81 75 -79
rect 77 -81 82 -79
rect 84 -81 95 -79
rect 73 -83 95 -81
rect 99 -79 105 -77
rect 99 -81 101 -79
rect 103 -81 105 -79
rect 99 -83 105 -81
rect 113 -80 115 -67
rect 123 -70 125 -67
rect 119 -72 125 -70
rect 119 -74 121 -72
rect 123 -74 125 -72
rect 119 -76 125 -74
rect 113 -82 119 -80
rect 14 -86 16 -83
rect 27 -86 29 -83
rect 34 -86 36 -83
rect 55 -86 57 -83
rect 65 -86 67 -83
rect 75 -86 77 -83
rect 93 -86 95 -83
rect 100 -86 102 -83
rect 113 -84 115 -82
rect 117 -84 119 -82
rect 110 -86 119 -84
rect 14 -118 16 -114
rect 110 -89 112 -86
rect 123 -89 125 -76
rect 151 -77 153 -68
rect 189 -60 191 -55
rect 199 -60 201 -55
rect 209 -57 211 -52
rect 219 -54 221 -50
rect 294 -54 296 -50
rect 305 -54 307 -50
rect 312 -54 314 -50
rect 253 -60 255 -55
rect 162 -77 164 -74
rect 169 -77 171 -74
rect 189 -77 191 -74
rect 199 -77 201 -74
rect 149 -79 155 -77
rect 149 -81 151 -79
rect 153 -81 155 -79
rect 149 -83 155 -81
rect 159 -79 165 -77
rect 159 -81 161 -79
rect 163 -81 165 -79
rect 159 -83 165 -81
rect 169 -79 191 -77
rect 169 -81 171 -79
rect 173 -81 178 -79
rect 180 -81 191 -79
rect 169 -83 191 -81
rect 195 -79 201 -77
rect 195 -81 197 -79
rect 199 -81 201 -79
rect 195 -83 201 -81
rect 209 -80 211 -67
rect 219 -70 221 -67
rect 215 -72 221 -70
rect 215 -74 217 -72
rect 219 -74 221 -72
rect 263 -61 265 -56
rect 273 -63 275 -59
rect 215 -76 221 -74
rect 209 -82 215 -80
rect 151 -86 153 -83
rect 161 -86 163 -83
rect 171 -86 173 -83
rect 189 -86 191 -83
rect 196 -86 198 -83
rect 209 -84 211 -82
rect 213 -84 215 -82
rect 206 -86 215 -84
rect 110 -107 112 -102
rect 27 -118 29 -114
rect 34 -118 36 -114
rect 55 -118 57 -114
rect 65 -118 67 -114
rect 75 -118 77 -114
rect 93 -116 95 -111
rect 100 -116 102 -111
rect 206 -89 208 -86
rect 219 -89 221 -76
rect 253 -77 255 -74
rect 263 -77 265 -69
rect 273 -77 275 -71
rect 294 -77 296 -68
rect 332 -60 334 -55
rect 342 -60 344 -55
rect 352 -57 354 -52
rect 362 -54 364 -50
rect 390 -54 392 -50
rect 401 -54 403 -50
rect 408 -54 410 -50
rect 305 -77 307 -74
rect 312 -77 314 -74
rect 332 -77 334 -74
rect 342 -77 344 -74
rect 253 -79 259 -77
rect 253 -81 255 -79
rect 257 -81 259 -79
rect 253 -83 259 -81
rect 263 -79 269 -77
rect 263 -81 265 -79
rect 267 -81 269 -79
rect 263 -83 269 -81
rect 273 -79 282 -77
rect 273 -81 278 -79
rect 280 -81 282 -79
rect 273 -83 282 -81
rect 292 -79 298 -77
rect 292 -81 294 -79
rect 296 -81 298 -79
rect 292 -83 298 -81
rect 302 -79 308 -77
rect 302 -81 304 -79
rect 306 -81 308 -79
rect 302 -83 308 -81
rect 312 -79 334 -77
rect 312 -81 314 -79
rect 316 -81 321 -79
rect 323 -81 334 -79
rect 312 -83 334 -81
rect 338 -79 344 -77
rect 338 -81 340 -79
rect 342 -81 344 -79
rect 338 -83 344 -81
rect 352 -80 354 -67
rect 362 -70 364 -67
rect 358 -72 364 -70
rect 358 -74 360 -72
rect 362 -74 364 -72
rect 358 -76 364 -74
rect 352 -82 358 -80
rect 253 -86 255 -83
rect 266 -86 268 -83
rect 273 -86 275 -83
rect 294 -86 296 -83
rect 304 -86 306 -83
rect 314 -86 316 -83
rect 332 -86 334 -83
rect 339 -86 341 -83
rect 352 -84 354 -82
rect 356 -84 358 -82
rect 349 -86 358 -84
rect 206 -107 208 -102
rect 123 -118 125 -114
rect 151 -118 153 -114
rect 161 -118 163 -114
rect 171 -118 173 -114
rect 189 -116 191 -111
rect 196 -116 198 -111
rect 219 -118 221 -114
rect 253 -118 255 -114
rect 349 -89 351 -86
rect 362 -89 364 -76
rect 390 -77 392 -68
rect 428 -60 430 -55
rect 438 -60 440 -55
rect 448 -57 450 -52
rect 458 -54 460 -50
rect 511 -52 530 -50
rect 511 -60 513 -52
rect 521 -60 523 -56
rect 528 -60 530 -52
rect 538 -60 540 -55
rect 545 -60 547 -55
rect 555 -60 557 -55
rect 401 -77 403 -74
rect 408 -77 410 -74
rect 428 -77 430 -74
rect 438 -77 440 -74
rect 388 -79 394 -77
rect 388 -81 390 -79
rect 392 -81 394 -79
rect 388 -83 394 -81
rect 398 -79 404 -77
rect 398 -81 400 -79
rect 402 -81 404 -79
rect 398 -83 404 -81
rect 408 -79 430 -77
rect 408 -81 410 -79
rect 412 -81 417 -79
rect 419 -81 430 -79
rect 408 -83 430 -81
rect 434 -79 440 -77
rect 434 -81 436 -79
rect 438 -81 440 -79
rect 434 -83 440 -81
rect 448 -80 450 -67
rect 458 -70 460 -67
rect 454 -72 460 -70
rect 454 -74 456 -72
rect 458 -74 460 -72
rect 454 -76 460 -74
rect 448 -82 454 -80
rect 390 -86 392 -83
rect 400 -86 402 -83
rect 410 -86 412 -83
rect 428 -86 430 -83
rect 435 -86 437 -83
rect 448 -84 450 -82
rect 452 -84 454 -82
rect 445 -86 454 -84
rect 349 -107 351 -102
rect 266 -118 268 -114
rect 273 -118 275 -114
rect 294 -118 296 -114
rect 304 -118 306 -114
rect 314 -118 316 -114
rect 332 -116 334 -111
rect 339 -116 341 -111
rect 445 -89 447 -86
rect 458 -89 460 -76
rect 511 -86 513 -66
rect 521 -77 523 -66
rect 517 -79 523 -77
rect 517 -81 519 -79
rect 521 -81 523 -79
rect 528 -79 530 -66
rect 538 -69 540 -66
rect 534 -71 540 -69
rect 534 -73 536 -71
rect 538 -73 540 -71
rect 534 -75 540 -73
rect 545 -79 547 -66
rect 555 -69 557 -66
rect 552 -71 558 -69
rect 552 -73 554 -71
rect 556 -73 558 -71
rect 552 -75 558 -73
rect 528 -81 540 -79
rect 517 -83 523 -81
rect 445 -107 447 -102
rect 362 -118 364 -114
rect 390 -118 392 -114
rect 400 -118 402 -114
rect 410 -118 412 -114
rect 428 -116 430 -111
rect 435 -116 437 -111
rect 511 -95 513 -92
rect 504 -97 513 -95
rect 521 -94 523 -83
rect 527 -87 533 -85
rect 527 -89 529 -87
rect 531 -89 533 -87
rect 527 -91 533 -89
rect 528 -94 530 -91
rect 538 -94 540 -81
rect 544 -81 550 -79
rect 544 -83 546 -81
rect 548 -83 550 -81
rect 544 -85 550 -83
rect 545 -94 547 -85
rect 555 -94 557 -75
rect 504 -99 506 -97
rect 508 -99 510 -97
rect 504 -101 510 -99
rect 521 -111 523 -106
rect 528 -111 530 -106
rect 538 -111 540 -106
rect 545 -111 547 -106
rect 555 -111 557 -106
rect 458 -118 460 -114
<< ndif >>
rect 84 235 90 237
rect 84 233 86 235
rect 88 233 90 235
rect 11 226 19 228
rect 11 224 14 226
rect 16 224 19 226
rect 11 219 19 224
rect 11 217 14 219
rect 16 217 19 219
rect 11 214 19 217
rect 21 225 28 228
rect 21 223 24 225
rect 26 223 28 225
rect 21 218 28 223
rect 21 216 24 218
rect 26 216 28 218
rect 21 214 28 216
rect 44 226 52 228
rect 44 224 47 226
rect 49 224 52 226
rect 44 219 52 224
rect 44 217 47 219
rect 49 217 52 219
rect 44 214 52 217
rect 54 225 61 228
rect 54 223 57 225
rect 59 223 61 225
rect 54 218 61 223
rect 84 227 90 233
rect 107 235 113 237
rect 107 233 109 235
rect 111 233 113 235
rect 107 231 113 233
rect 107 227 111 231
rect 84 221 93 227
rect 95 225 103 227
rect 95 223 98 225
rect 100 223 103 225
rect 95 221 103 223
rect 105 225 111 227
rect 146 225 153 228
rect 105 221 113 225
rect 54 216 57 218
rect 59 216 61 218
rect 54 214 61 216
rect 107 219 113 221
rect 115 223 123 225
rect 115 221 118 223
rect 120 221 123 223
rect 115 219 123 221
rect 125 223 132 225
rect 125 221 128 223
rect 130 221 132 223
rect 125 219 132 221
rect 146 223 148 225
rect 150 223 153 225
rect 146 218 153 223
rect 146 216 148 218
rect 150 216 153 218
rect 146 214 153 216
rect 155 226 163 228
rect 155 224 158 226
rect 160 224 163 226
rect 155 219 163 224
rect 155 217 158 219
rect 160 217 163 219
rect 155 214 163 217
rect 181 226 189 228
rect 181 224 184 226
rect 186 224 189 226
rect 181 219 189 224
rect 181 217 184 219
rect 186 217 189 219
rect 181 214 189 217
rect 191 225 198 228
rect 191 223 194 225
rect 196 223 198 225
rect 191 218 198 223
rect 212 226 219 228
rect 212 224 214 226
rect 216 224 219 226
rect 212 222 219 224
rect 221 226 229 228
rect 221 224 224 226
rect 226 224 229 226
rect 221 222 229 224
rect 231 222 236 228
rect 238 226 246 228
rect 238 224 241 226
rect 243 224 246 226
rect 238 222 246 224
rect 248 222 253 228
rect 255 226 263 228
rect 255 224 258 226
rect 260 224 263 226
rect 255 222 263 224
rect 265 226 272 228
rect 265 224 268 226
rect 270 224 272 226
rect 297 225 302 231
rect 265 222 272 224
rect 284 222 292 225
rect 191 216 194 218
rect 196 216 198 218
rect 191 214 198 216
rect 284 220 287 222
rect 289 220 292 222
rect 284 214 292 220
rect 294 218 302 225
rect 294 216 297 218
rect 299 216 302 218
rect 294 214 302 216
rect 304 229 311 231
rect 304 227 307 229
rect 309 227 311 229
rect 304 214 311 227
rect 322 226 329 228
rect 322 224 324 226
rect 326 224 329 226
rect 322 222 329 224
rect 331 226 339 228
rect 331 224 334 226
rect 336 224 339 226
rect 331 222 339 224
rect 341 222 346 228
rect 348 226 356 228
rect 348 224 351 226
rect 353 224 356 226
rect 348 222 356 224
rect 358 222 363 228
rect 365 226 373 228
rect 365 224 368 226
rect 370 224 373 226
rect 365 222 373 224
rect 375 226 382 228
rect 375 224 378 226
rect 380 224 382 226
rect 375 222 382 224
rect 390 226 397 229
rect 390 224 392 226
rect 394 224 397 226
rect 390 219 397 224
rect 390 217 392 219
rect 394 217 397 219
rect 390 215 397 217
rect 399 227 407 229
rect 399 225 402 227
rect 404 225 407 227
rect 399 215 407 225
rect 409 225 417 229
rect 409 223 412 225
rect 414 223 417 225
rect 409 215 417 223
rect 419 227 426 229
rect 419 225 422 227
rect 424 225 426 227
rect 419 219 426 225
rect 419 217 422 219
rect 424 217 426 219
rect 419 215 426 217
rect 442 226 449 229
rect 442 224 444 226
rect 446 224 449 226
rect 442 219 449 224
rect 442 217 444 219
rect 446 217 449 219
rect 442 215 449 217
rect 451 227 459 229
rect 451 225 454 227
rect 456 225 459 227
rect 451 215 459 225
rect 461 225 469 229
rect 461 223 464 225
rect 466 223 469 225
rect 461 215 469 223
rect 471 227 478 229
rect 471 225 474 227
rect 476 225 478 227
rect 471 219 478 225
rect 471 217 474 219
rect 476 217 478 219
rect 471 215 478 217
rect 484 226 491 229
rect 484 224 486 226
rect 488 224 491 226
rect 484 219 491 224
rect 484 217 486 219
rect 488 217 491 219
rect 484 215 491 217
rect 493 227 501 229
rect 493 225 496 227
rect 498 225 501 227
rect 493 215 501 225
rect 503 225 511 229
rect 503 223 506 225
rect 508 223 511 225
rect 503 215 511 223
rect 513 227 520 229
rect 513 225 516 227
rect 518 225 520 227
rect 513 219 520 225
rect 513 217 516 219
rect 518 217 520 219
rect 513 215 520 217
rect 528 226 535 229
rect 528 224 530 226
rect 532 224 535 226
rect 528 219 535 224
rect 528 217 530 219
rect 532 217 535 219
rect 528 215 535 217
rect 537 227 545 229
rect 537 225 540 227
rect 542 225 545 227
rect 537 215 545 225
rect 547 225 555 229
rect 547 223 550 225
rect 552 223 555 225
rect 547 215 555 223
rect 557 227 564 229
rect 557 225 560 227
rect 562 225 564 227
rect 557 219 564 225
rect 557 217 560 219
rect 562 217 564 219
rect 557 215 564 217
rect 29 115 34 122
rect 7 113 14 115
rect 7 111 9 113
rect 11 111 14 113
rect 7 109 14 111
rect 9 102 14 109
rect 16 109 24 115
rect 16 107 19 109
rect 21 107 24 109
rect 16 105 24 107
rect 26 112 34 115
rect 26 110 29 112
rect 31 110 34 112
rect 26 108 34 110
rect 36 120 44 122
rect 36 118 39 120
rect 41 118 44 120
rect 36 108 44 118
rect 46 120 53 122
rect 46 118 49 120
rect 51 118 53 120
rect 46 113 53 118
rect 59 115 64 122
rect 46 111 49 113
rect 51 111 53 113
rect 46 108 53 111
rect 57 113 64 115
rect 57 111 59 113
rect 61 111 64 113
rect 57 109 64 111
rect 26 105 31 108
rect 16 102 21 105
rect 59 102 64 109
rect 66 102 71 122
rect 73 116 80 122
rect 73 106 82 116
rect 73 104 76 106
rect 78 104 82 106
rect 73 102 82 104
rect 84 113 91 116
rect 125 115 130 122
rect 84 111 87 113
rect 89 111 91 113
rect 84 109 91 111
rect 103 113 110 115
rect 103 111 105 113
rect 107 111 110 113
rect 103 109 110 111
rect 84 102 89 109
rect 105 102 110 109
rect 112 109 120 115
rect 112 107 115 109
rect 117 107 120 109
rect 112 105 120 107
rect 122 112 130 115
rect 122 110 125 112
rect 127 110 130 112
rect 122 108 130 110
rect 132 120 140 122
rect 132 118 135 120
rect 137 118 140 120
rect 132 108 140 118
rect 142 120 149 122
rect 142 118 145 120
rect 147 118 149 120
rect 142 113 149 118
rect 155 115 160 122
rect 142 111 145 113
rect 147 111 149 113
rect 142 108 149 111
rect 153 113 160 115
rect 153 111 155 113
rect 157 111 160 113
rect 153 109 160 111
rect 122 105 127 108
rect 112 102 117 105
rect 155 102 160 109
rect 162 102 167 122
rect 169 116 176 122
rect 169 106 178 116
rect 169 104 172 106
rect 174 104 178 106
rect 169 102 178 104
rect 180 113 187 116
rect 180 111 183 113
rect 185 111 187 113
rect 192 115 199 119
rect 192 113 194 115
rect 196 113 199 115
rect 192 111 199 113
rect 201 117 206 119
rect 214 117 219 122
rect 201 115 209 117
rect 201 113 204 115
rect 206 113 209 115
rect 201 111 209 113
rect 180 109 187 111
rect 180 102 185 109
rect 204 109 209 111
rect 211 113 219 117
rect 211 111 214 113
rect 216 111 219 113
rect 211 109 219 111
rect 214 108 219 109
rect 221 120 228 122
rect 221 118 224 120
rect 226 118 228 120
rect 221 113 228 118
rect 269 115 274 122
rect 221 111 224 113
rect 226 111 228 113
rect 221 108 228 111
rect 247 113 254 115
rect 247 111 249 113
rect 251 111 254 113
rect 247 109 254 111
rect 249 102 254 109
rect 256 109 264 115
rect 256 107 259 109
rect 261 107 264 109
rect 256 105 264 107
rect 266 112 274 115
rect 266 110 269 112
rect 271 110 274 112
rect 266 108 274 110
rect 276 120 284 122
rect 276 118 279 120
rect 281 118 284 120
rect 276 108 284 118
rect 286 120 293 122
rect 286 118 289 120
rect 291 118 293 120
rect 286 113 293 118
rect 299 115 304 122
rect 286 111 289 113
rect 291 111 293 113
rect 286 108 293 111
rect 297 113 304 115
rect 297 111 299 113
rect 301 111 304 113
rect 297 109 304 111
rect 266 105 271 108
rect 256 102 261 105
rect 299 102 304 109
rect 306 102 311 122
rect 313 116 320 122
rect 313 106 322 116
rect 313 104 316 106
rect 318 104 322 106
rect 313 102 322 104
rect 324 113 331 116
rect 365 115 370 122
rect 324 111 327 113
rect 329 111 331 113
rect 324 109 331 111
rect 343 113 350 115
rect 343 111 345 113
rect 347 111 350 113
rect 343 109 350 111
rect 324 102 329 109
rect 345 102 350 109
rect 352 109 360 115
rect 352 107 355 109
rect 357 107 360 109
rect 352 105 360 107
rect 362 112 370 115
rect 362 110 365 112
rect 367 110 370 112
rect 362 108 370 110
rect 372 120 380 122
rect 372 118 375 120
rect 377 118 380 120
rect 372 108 380 118
rect 382 120 389 122
rect 382 118 385 120
rect 387 118 389 120
rect 382 113 389 118
rect 395 115 400 122
rect 382 111 385 113
rect 387 111 389 113
rect 382 108 389 111
rect 393 113 400 115
rect 393 111 395 113
rect 397 111 400 113
rect 393 109 400 111
rect 362 105 367 108
rect 352 102 357 105
rect 395 102 400 109
rect 402 102 407 122
rect 409 116 416 122
rect 409 106 418 116
rect 409 104 412 106
rect 414 104 418 106
rect 409 102 418 104
rect 420 113 427 116
rect 420 111 423 113
rect 425 111 427 113
rect 432 115 439 119
rect 432 113 434 115
rect 436 113 439 115
rect 432 111 439 113
rect 441 117 446 119
rect 454 117 459 122
rect 441 115 449 117
rect 441 113 444 115
rect 446 113 449 115
rect 441 111 449 113
rect 420 109 427 111
rect 420 102 425 109
rect 444 109 449 111
rect 451 113 459 117
rect 451 111 454 113
rect 456 111 459 113
rect 451 109 459 111
rect 454 108 459 109
rect 461 120 468 122
rect 461 118 464 120
rect 466 118 468 120
rect 461 113 468 118
rect 461 111 464 113
rect 466 111 468 113
rect 461 108 468 111
rect 504 112 511 114
rect 504 110 506 112
rect 508 110 511 112
rect 504 108 511 110
rect 513 112 521 114
rect 513 110 516 112
rect 518 110 521 112
rect 513 108 521 110
rect 523 108 528 114
rect 530 112 538 114
rect 530 110 533 112
rect 535 110 538 112
rect 530 108 538 110
rect 540 108 545 114
rect 547 112 555 114
rect 547 110 550 112
rect 552 110 555 112
rect 547 108 555 110
rect 557 112 564 114
rect 557 110 560 112
rect 562 110 564 112
rect 557 108 564 110
rect 7 81 14 84
rect 7 79 9 81
rect 11 79 14 81
rect 7 74 14 79
rect 7 72 9 74
rect 11 72 14 74
rect 7 70 14 72
rect 16 83 21 84
rect 16 81 24 83
rect 16 79 19 81
rect 21 79 24 81
rect 16 75 24 79
rect 26 81 31 83
rect 50 83 55 90
rect 48 81 55 83
rect 26 79 34 81
rect 26 77 29 79
rect 31 77 34 79
rect 26 75 34 77
rect 16 70 21 75
rect 29 73 34 75
rect 36 79 43 81
rect 36 77 39 79
rect 41 77 43 79
rect 36 73 43 77
rect 48 79 50 81
rect 52 79 55 81
rect 48 76 55 79
rect 57 88 66 90
rect 57 86 61 88
rect 63 86 66 88
rect 57 76 66 86
rect 59 70 66 76
rect 68 70 73 90
rect 75 83 80 90
rect 118 87 123 90
rect 108 84 113 87
rect 75 81 82 83
rect 75 79 78 81
rect 80 79 82 81
rect 75 77 82 79
rect 86 81 93 84
rect 86 79 88 81
rect 90 79 93 81
rect 75 70 80 77
rect 86 74 93 79
rect 86 72 88 74
rect 90 72 93 74
rect 86 70 93 72
rect 95 74 103 84
rect 95 72 98 74
rect 100 72 103 74
rect 95 70 103 72
rect 105 82 113 84
rect 105 80 108 82
rect 110 80 113 82
rect 105 77 113 80
rect 115 85 123 87
rect 115 83 118 85
rect 120 83 123 85
rect 115 77 123 83
rect 125 83 130 90
rect 146 83 151 90
rect 125 81 132 83
rect 125 79 128 81
rect 130 79 132 81
rect 125 77 132 79
rect 144 81 151 83
rect 144 79 146 81
rect 148 79 151 81
rect 105 70 110 77
rect 144 76 151 79
rect 153 88 162 90
rect 153 86 157 88
rect 159 86 162 88
rect 153 76 162 86
rect 155 70 162 76
rect 164 70 169 90
rect 171 83 176 90
rect 214 87 219 90
rect 204 84 209 87
rect 171 81 178 83
rect 171 79 174 81
rect 176 79 178 81
rect 171 77 178 79
rect 182 81 189 84
rect 182 79 184 81
rect 186 79 189 81
rect 171 70 176 77
rect 182 74 189 79
rect 182 72 184 74
rect 186 72 189 74
rect 182 70 189 72
rect 191 74 199 84
rect 191 72 194 74
rect 196 72 199 74
rect 191 70 199 72
rect 201 82 209 84
rect 201 80 204 82
rect 206 80 209 82
rect 201 77 209 80
rect 211 85 219 87
rect 211 83 214 85
rect 216 83 219 85
rect 211 77 219 83
rect 221 83 226 90
rect 221 81 228 83
rect 221 79 224 81
rect 226 79 228 81
rect 221 77 228 79
rect 246 81 253 84
rect 246 79 248 81
rect 250 79 253 81
rect 201 70 206 77
rect 246 74 253 79
rect 246 72 248 74
rect 250 72 253 74
rect 246 70 253 72
rect 255 83 260 84
rect 255 81 263 83
rect 255 79 258 81
rect 260 79 263 81
rect 255 75 263 79
rect 265 81 270 83
rect 289 83 294 90
rect 287 81 294 83
rect 265 79 273 81
rect 265 77 268 79
rect 270 77 273 79
rect 265 75 273 77
rect 255 70 260 75
rect 268 73 273 75
rect 275 79 282 81
rect 275 77 278 79
rect 280 77 282 79
rect 275 73 282 77
rect 287 79 289 81
rect 291 79 294 81
rect 287 76 294 79
rect 296 88 305 90
rect 296 86 300 88
rect 302 86 305 88
rect 296 76 305 86
rect 298 70 305 76
rect 307 70 312 90
rect 314 83 319 90
rect 357 87 362 90
rect 347 84 352 87
rect 314 81 321 83
rect 314 79 317 81
rect 319 79 321 81
rect 314 77 321 79
rect 325 81 332 84
rect 325 79 327 81
rect 329 79 332 81
rect 314 70 319 77
rect 325 74 332 79
rect 325 72 327 74
rect 329 72 332 74
rect 325 70 332 72
rect 334 74 342 84
rect 334 72 337 74
rect 339 72 342 74
rect 334 70 342 72
rect 344 82 352 84
rect 344 80 347 82
rect 349 80 352 82
rect 344 77 352 80
rect 354 85 362 87
rect 354 83 357 85
rect 359 83 362 85
rect 354 77 362 83
rect 364 83 369 90
rect 385 83 390 90
rect 364 81 371 83
rect 364 79 367 81
rect 369 79 371 81
rect 364 77 371 79
rect 383 81 390 83
rect 383 79 385 81
rect 387 79 390 81
rect 344 70 349 77
rect 383 76 390 79
rect 392 88 401 90
rect 392 86 396 88
rect 398 86 401 88
rect 392 76 401 86
rect 394 70 401 76
rect 403 70 408 90
rect 410 83 415 90
rect 453 87 458 90
rect 443 84 448 87
rect 410 81 417 83
rect 410 79 413 81
rect 415 79 417 81
rect 410 77 417 79
rect 421 81 428 84
rect 421 79 423 81
rect 425 79 428 81
rect 410 70 415 77
rect 421 74 428 79
rect 421 72 423 74
rect 425 72 428 74
rect 421 70 428 72
rect 430 74 438 84
rect 430 72 433 74
rect 435 72 438 74
rect 430 70 438 72
rect 440 82 448 84
rect 440 80 443 82
rect 445 80 448 82
rect 440 77 448 80
rect 450 85 458 87
rect 450 83 453 85
rect 455 83 458 85
rect 450 77 458 83
rect 460 83 465 90
rect 460 81 467 83
rect 460 79 463 81
rect 465 79 467 81
rect 460 77 467 79
rect 504 82 511 84
rect 504 80 506 82
rect 508 80 511 82
rect 504 78 511 80
rect 513 82 521 84
rect 513 80 516 82
rect 518 80 521 82
rect 513 78 521 80
rect 523 78 528 84
rect 530 82 538 84
rect 530 80 533 82
rect 535 80 538 82
rect 530 78 538 80
rect 540 78 545 84
rect 547 82 555 84
rect 547 80 550 82
rect 552 80 555 82
rect 547 78 555 80
rect 557 82 564 84
rect 557 80 560 82
rect 562 80 564 82
rect 557 78 564 80
rect 440 70 445 77
rect 29 -29 34 -22
rect 7 -31 14 -29
rect 7 -33 9 -31
rect 11 -33 14 -31
rect 7 -35 14 -33
rect 9 -42 14 -35
rect 16 -35 24 -29
rect 16 -37 19 -35
rect 21 -37 24 -35
rect 16 -39 24 -37
rect 26 -32 34 -29
rect 26 -34 29 -32
rect 31 -34 34 -32
rect 26 -36 34 -34
rect 36 -24 44 -22
rect 36 -26 39 -24
rect 41 -26 44 -24
rect 36 -36 44 -26
rect 46 -24 53 -22
rect 46 -26 49 -24
rect 51 -26 53 -24
rect 46 -31 53 -26
rect 59 -29 64 -22
rect 46 -33 49 -31
rect 51 -33 53 -31
rect 46 -36 53 -33
rect 57 -31 64 -29
rect 57 -33 59 -31
rect 61 -33 64 -31
rect 57 -35 64 -33
rect 26 -39 31 -36
rect 16 -42 21 -39
rect 59 -42 64 -35
rect 66 -42 71 -22
rect 73 -28 80 -22
rect 73 -38 82 -28
rect 73 -40 76 -38
rect 78 -40 82 -38
rect 73 -42 82 -40
rect 84 -31 91 -28
rect 125 -29 130 -22
rect 84 -33 87 -31
rect 89 -33 91 -31
rect 84 -35 91 -33
rect 103 -31 110 -29
rect 103 -33 105 -31
rect 107 -33 110 -31
rect 103 -35 110 -33
rect 84 -42 89 -35
rect 105 -42 110 -35
rect 112 -35 120 -29
rect 112 -37 115 -35
rect 117 -37 120 -35
rect 112 -39 120 -37
rect 122 -32 130 -29
rect 122 -34 125 -32
rect 127 -34 130 -32
rect 122 -36 130 -34
rect 132 -24 140 -22
rect 132 -26 135 -24
rect 137 -26 140 -24
rect 132 -36 140 -26
rect 142 -24 149 -22
rect 142 -26 145 -24
rect 147 -26 149 -24
rect 142 -31 149 -26
rect 155 -29 160 -22
rect 142 -33 145 -31
rect 147 -33 149 -31
rect 142 -36 149 -33
rect 153 -31 160 -29
rect 153 -33 155 -31
rect 157 -33 160 -31
rect 153 -35 160 -33
rect 122 -39 127 -36
rect 112 -42 117 -39
rect 155 -42 160 -35
rect 162 -42 167 -22
rect 169 -28 176 -22
rect 169 -38 178 -28
rect 169 -40 172 -38
rect 174 -40 178 -38
rect 169 -42 178 -40
rect 180 -31 187 -28
rect 180 -33 183 -31
rect 185 -33 187 -31
rect 192 -29 199 -25
rect 192 -31 194 -29
rect 196 -31 199 -29
rect 192 -33 199 -31
rect 201 -27 206 -25
rect 214 -27 219 -22
rect 201 -29 209 -27
rect 201 -31 204 -29
rect 206 -31 209 -29
rect 201 -33 209 -31
rect 180 -35 187 -33
rect 180 -42 185 -35
rect 204 -35 209 -33
rect 211 -31 219 -27
rect 211 -33 214 -31
rect 216 -33 219 -31
rect 211 -35 219 -33
rect 214 -36 219 -35
rect 221 -24 228 -22
rect 221 -26 224 -24
rect 226 -26 228 -24
rect 221 -31 228 -26
rect 269 -29 274 -22
rect 221 -33 224 -31
rect 226 -33 228 -31
rect 221 -36 228 -33
rect 247 -31 254 -29
rect 247 -33 249 -31
rect 251 -33 254 -31
rect 247 -35 254 -33
rect 249 -42 254 -35
rect 256 -35 264 -29
rect 256 -37 259 -35
rect 261 -37 264 -35
rect 256 -39 264 -37
rect 266 -32 274 -29
rect 266 -34 269 -32
rect 271 -34 274 -32
rect 266 -36 274 -34
rect 276 -24 284 -22
rect 276 -26 279 -24
rect 281 -26 284 -24
rect 276 -36 284 -26
rect 286 -24 293 -22
rect 286 -26 289 -24
rect 291 -26 293 -24
rect 286 -31 293 -26
rect 299 -29 304 -22
rect 286 -33 289 -31
rect 291 -33 293 -31
rect 286 -36 293 -33
rect 297 -31 304 -29
rect 297 -33 299 -31
rect 301 -33 304 -31
rect 297 -35 304 -33
rect 266 -39 271 -36
rect 256 -42 261 -39
rect 299 -42 304 -35
rect 306 -42 311 -22
rect 313 -28 320 -22
rect 313 -38 322 -28
rect 313 -40 316 -38
rect 318 -40 322 -38
rect 313 -42 322 -40
rect 324 -31 331 -28
rect 365 -29 370 -22
rect 324 -33 327 -31
rect 329 -33 331 -31
rect 324 -35 331 -33
rect 343 -31 350 -29
rect 343 -33 345 -31
rect 347 -33 350 -31
rect 343 -35 350 -33
rect 324 -42 329 -35
rect 345 -42 350 -35
rect 352 -35 360 -29
rect 352 -37 355 -35
rect 357 -37 360 -35
rect 352 -39 360 -37
rect 362 -32 370 -29
rect 362 -34 365 -32
rect 367 -34 370 -32
rect 362 -36 370 -34
rect 372 -24 380 -22
rect 372 -26 375 -24
rect 377 -26 380 -24
rect 372 -36 380 -26
rect 382 -24 389 -22
rect 382 -26 385 -24
rect 387 -26 389 -24
rect 382 -31 389 -26
rect 395 -29 400 -22
rect 382 -33 385 -31
rect 387 -33 389 -31
rect 382 -36 389 -33
rect 393 -31 400 -29
rect 393 -33 395 -31
rect 397 -33 400 -31
rect 393 -35 400 -33
rect 362 -39 367 -36
rect 352 -42 357 -39
rect 395 -42 400 -35
rect 402 -42 407 -22
rect 409 -28 416 -22
rect 409 -38 418 -28
rect 409 -40 412 -38
rect 414 -40 418 -38
rect 409 -42 418 -40
rect 420 -31 427 -28
rect 420 -33 423 -31
rect 425 -33 427 -31
rect 432 -29 439 -25
rect 432 -31 434 -29
rect 436 -31 439 -29
rect 432 -33 439 -31
rect 441 -27 446 -25
rect 454 -27 459 -22
rect 441 -29 449 -27
rect 441 -31 444 -29
rect 446 -31 449 -29
rect 441 -33 449 -31
rect 420 -35 427 -33
rect 420 -42 425 -35
rect 444 -35 449 -33
rect 451 -31 459 -27
rect 451 -33 454 -31
rect 456 -33 459 -31
rect 451 -35 459 -33
rect 454 -36 459 -35
rect 461 -24 468 -22
rect 461 -26 464 -24
rect 466 -26 468 -24
rect 461 -31 468 -26
rect 461 -33 464 -31
rect 466 -33 468 -31
rect 461 -36 468 -33
rect 504 -32 511 -30
rect 504 -34 506 -32
rect 508 -34 511 -32
rect 504 -36 511 -34
rect 513 -32 521 -30
rect 513 -34 516 -32
rect 518 -34 521 -32
rect 513 -36 521 -34
rect 523 -36 528 -30
rect 530 -32 538 -30
rect 530 -34 533 -32
rect 535 -34 538 -32
rect 530 -36 538 -34
rect 540 -36 545 -30
rect 547 -32 555 -30
rect 547 -34 550 -32
rect 552 -34 555 -32
rect 547 -36 555 -34
rect 557 -32 564 -30
rect 557 -34 560 -32
rect 562 -34 564 -32
rect 557 -36 564 -34
rect 7 -63 14 -60
rect 7 -65 9 -63
rect 11 -65 14 -63
rect 7 -70 14 -65
rect 7 -72 9 -70
rect 11 -72 14 -70
rect 7 -74 14 -72
rect 16 -61 21 -60
rect 16 -63 24 -61
rect 16 -65 19 -63
rect 21 -65 24 -63
rect 16 -69 24 -65
rect 26 -63 31 -61
rect 50 -61 55 -54
rect 48 -63 55 -61
rect 26 -65 34 -63
rect 26 -67 29 -65
rect 31 -67 34 -65
rect 26 -69 34 -67
rect 16 -74 21 -69
rect 29 -71 34 -69
rect 36 -65 43 -63
rect 36 -67 39 -65
rect 41 -67 43 -65
rect 36 -71 43 -67
rect 48 -65 50 -63
rect 52 -65 55 -63
rect 48 -68 55 -65
rect 57 -56 66 -54
rect 57 -58 61 -56
rect 63 -58 66 -56
rect 57 -68 66 -58
rect 59 -74 66 -68
rect 68 -74 73 -54
rect 75 -61 80 -54
rect 118 -57 123 -54
rect 108 -60 113 -57
rect 75 -63 82 -61
rect 75 -65 78 -63
rect 80 -65 82 -63
rect 75 -67 82 -65
rect 86 -63 93 -60
rect 86 -65 88 -63
rect 90 -65 93 -63
rect 75 -74 80 -67
rect 86 -70 93 -65
rect 86 -72 88 -70
rect 90 -72 93 -70
rect 86 -74 93 -72
rect 95 -70 103 -60
rect 95 -72 98 -70
rect 100 -72 103 -70
rect 95 -74 103 -72
rect 105 -62 113 -60
rect 105 -64 108 -62
rect 110 -64 113 -62
rect 105 -67 113 -64
rect 115 -59 123 -57
rect 115 -61 118 -59
rect 120 -61 123 -59
rect 115 -67 123 -61
rect 125 -61 130 -54
rect 146 -61 151 -54
rect 125 -63 132 -61
rect 125 -65 128 -63
rect 130 -65 132 -63
rect 125 -67 132 -65
rect 144 -63 151 -61
rect 144 -65 146 -63
rect 148 -65 151 -63
rect 105 -74 110 -67
rect 144 -68 151 -65
rect 153 -56 162 -54
rect 153 -58 157 -56
rect 159 -58 162 -56
rect 153 -68 162 -58
rect 155 -74 162 -68
rect 164 -74 169 -54
rect 171 -61 176 -54
rect 214 -57 219 -54
rect 204 -60 209 -57
rect 171 -63 178 -61
rect 171 -65 174 -63
rect 176 -65 178 -63
rect 171 -67 178 -65
rect 182 -63 189 -60
rect 182 -65 184 -63
rect 186 -65 189 -63
rect 171 -74 176 -67
rect 182 -70 189 -65
rect 182 -72 184 -70
rect 186 -72 189 -70
rect 182 -74 189 -72
rect 191 -70 199 -60
rect 191 -72 194 -70
rect 196 -72 199 -70
rect 191 -74 199 -72
rect 201 -62 209 -60
rect 201 -64 204 -62
rect 206 -64 209 -62
rect 201 -67 209 -64
rect 211 -59 219 -57
rect 211 -61 214 -59
rect 216 -61 219 -59
rect 211 -67 219 -61
rect 221 -61 226 -54
rect 221 -63 228 -61
rect 221 -65 224 -63
rect 226 -65 228 -63
rect 221 -67 228 -65
rect 246 -63 253 -60
rect 246 -65 248 -63
rect 250 -65 253 -63
rect 201 -74 206 -67
rect 246 -70 253 -65
rect 246 -72 248 -70
rect 250 -72 253 -70
rect 246 -74 253 -72
rect 255 -61 260 -60
rect 255 -63 263 -61
rect 255 -65 258 -63
rect 260 -65 263 -63
rect 255 -69 263 -65
rect 265 -63 270 -61
rect 289 -61 294 -54
rect 287 -63 294 -61
rect 265 -65 273 -63
rect 265 -67 268 -65
rect 270 -67 273 -65
rect 265 -69 273 -67
rect 255 -74 260 -69
rect 268 -71 273 -69
rect 275 -65 282 -63
rect 275 -67 278 -65
rect 280 -67 282 -65
rect 275 -71 282 -67
rect 287 -65 289 -63
rect 291 -65 294 -63
rect 287 -68 294 -65
rect 296 -56 305 -54
rect 296 -58 300 -56
rect 302 -58 305 -56
rect 296 -68 305 -58
rect 298 -74 305 -68
rect 307 -74 312 -54
rect 314 -61 319 -54
rect 357 -57 362 -54
rect 347 -60 352 -57
rect 314 -63 321 -61
rect 314 -65 317 -63
rect 319 -65 321 -63
rect 314 -67 321 -65
rect 325 -63 332 -60
rect 325 -65 327 -63
rect 329 -65 332 -63
rect 314 -74 319 -67
rect 325 -70 332 -65
rect 325 -72 327 -70
rect 329 -72 332 -70
rect 325 -74 332 -72
rect 334 -70 342 -60
rect 334 -72 337 -70
rect 339 -72 342 -70
rect 334 -74 342 -72
rect 344 -62 352 -60
rect 344 -64 347 -62
rect 349 -64 352 -62
rect 344 -67 352 -64
rect 354 -59 362 -57
rect 354 -61 357 -59
rect 359 -61 362 -59
rect 354 -67 362 -61
rect 364 -61 369 -54
rect 385 -61 390 -54
rect 364 -63 371 -61
rect 364 -65 367 -63
rect 369 -65 371 -63
rect 364 -67 371 -65
rect 383 -63 390 -61
rect 383 -65 385 -63
rect 387 -65 390 -63
rect 344 -74 349 -67
rect 383 -68 390 -65
rect 392 -56 401 -54
rect 392 -58 396 -56
rect 398 -58 401 -56
rect 392 -68 401 -58
rect 394 -74 401 -68
rect 403 -74 408 -54
rect 410 -61 415 -54
rect 453 -57 458 -54
rect 443 -60 448 -57
rect 410 -63 417 -61
rect 410 -65 413 -63
rect 415 -65 417 -63
rect 410 -67 417 -65
rect 421 -63 428 -60
rect 421 -65 423 -63
rect 425 -65 428 -63
rect 410 -74 415 -67
rect 421 -70 428 -65
rect 421 -72 423 -70
rect 425 -72 428 -70
rect 421 -74 428 -72
rect 430 -70 438 -60
rect 430 -72 433 -70
rect 435 -72 438 -70
rect 430 -74 438 -72
rect 440 -62 448 -60
rect 440 -64 443 -62
rect 445 -64 448 -62
rect 440 -67 448 -64
rect 450 -59 458 -57
rect 450 -61 453 -59
rect 455 -61 458 -59
rect 450 -67 458 -61
rect 460 -61 465 -54
rect 460 -63 467 -61
rect 460 -65 463 -63
rect 465 -65 467 -63
rect 460 -67 467 -65
rect 504 -62 511 -60
rect 504 -64 506 -62
rect 508 -64 511 -62
rect 504 -66 511 -64
rect 513 -62 521 -60
rect 513 -64 516 -62
rect 518 -64 521 -62
rect 513 -66 521 -64
rect 523 -66 528 -60
rect 530 -62 538 -60
rect 530 -64 533 -62
rect 535 -64 538 -62
rect 530 -66 538 -64
rect 540 -66 545 -60
rect 547 -62 555 -60
rect 547 -64 550 -62
rect 552 -64 555 -62
rect 547 -66 555 -64
rect 557 -62 564 -60
rect 557 -64 560 -62
rect 562 -64 564 -62
rect 557 -66 564 -64
rect 440 -74 445 -67
<< pdif >>
rect 11 185 19 202
rect 11 183 14 185
rect 16 183 19 185
rect 11 178 19 183
rect 11 176 14 178
rect 16 176 19 178
rect 11 174 19 176
rect 21 199 28 202
rect 21 197 24 199
rect 26 197 28 199
rect 21 192 28 197
rect 21 190 24 192
rect 26 190 28 192
rect 21 188 28 190
rect 21 174 26 188
rect 44 185 52 202
rect 44 183 47 185
rect 49 183 52 185
rect 44 178 52 183
rect 44 176 47 178
rect 49 176 52 178
rect 44 174 52 176
rect 54 199 61 202
rect 54 197 57 199
rect 59 197 61 199
rect 54 193 61 197
rect 146 199 153 202
rect 146 197 148 199
rect 150 197 153 199
rect 54 192 67 193
rect 54 190 57 192
rect 59 190 67 192
rect 54 189 67 190
rect 54 188 61 189
rect 54 174 59 188
rect 86 186 93 196
rect 86 184 88 186
rect 90 184 93 186
rect 86 178 93 184
rect 86 176 88 178
rect 90 176 93 178
rect 86 174 93 176
rect 95 174 100 196
rect 102 174 107 196
rect 109 174 114 196
rect 116 187 121 196
rect 146 192 153 197
rect 146 190 148 192
rect 150 190 153 192
rect 146 188 153 190
rect 116 185 123 187
rect 116 183 119 185
rect 121 183 123 185
rect 116 181 123 183
rect 116 174 121 181
rect 148 174 153 188
rect 155 185 163 202
rect 155 183 158 185
rect 160 183 163 185
rect 155 178 163 183
rect 155 176 158 178
rect 160 176 163 178
rect 155 174 163 176
rect 181 185 189 202
rect 181 183 184 185
rect 186 183 189 185
rect 181 178 189 183
rect 181 176 184 178
rect 186 176 189 178
rect 181 174 189 176
rect 191 199 198 202
rect 191 197 194 199
rect 196 197 198 199
rect 191 192 198 197
rect 212 200 219 202
rect 212 198 214 200
rect 216 198 219 200
rect 212 196 219 198
rect 221 196 227 202
rect 191 190 194 192
rect 196 190 198 192
rect 191 188 198 190
rect 223 194 227 196
rect 191 174 196 188
rect 223 188 229 194
rect 222 186 229 188
rect 222 184 224 186
rect 226 184 229 186
rect 222 182 229 184
rect 231 182 236 194
rect 238 192 246 194
rect 238 190 241 192
rect 243 190 246 192
rect 238 182 246 190
rect 248 182 253 194
rect 255 186 263 194
rect 255 184 258 186
rect 260 184 263 186
rect 255 182 263 184
rect 265 192 272 194
rect 265 190 268 192
rect 270 190 272 192
rect 265 188 272 190
rect 265 182 270 188
rect 284 185 292 202
rect 284 183 287 185
rect 289 183 292 185
rect 284 178 292 183
rect 284 176 287 178
rect 289 176 292 178
rect 284 174 292 176
rect 294 192 302 202
rect 294 190 297 192
rect 299 190 302 192
rect 294 185 302 190
rect 294 183 297 185
rect 299 183 302 185
rect 294 174 302 183
rect 304 185 311 202
rect 322 200 329 202
rect 322 198 324 200
rect 326 198 329 200
rect 322 196 329 198
rect 331 196 337 202
rect 333 194 337 196
rect 390 200 397 202
rect 390 198 392 200
rect 394 198 397 200
rect 333 188 339 194
rect 304 183 307 185
rect 309 183 311 185
rect 304 178 311 183
rect 332 186 339 188
rect 332 184 334 186
rect 336 184 339 186
rect 332 182 339 184
rect 341 182 346 194
rect 348 192 356 194
rect 348 190 351 192
rect 353 190 356 192
rect 348 182 356 190
rect 358 182 363 194
rect 365 186 373 194
rect 365 184 368 186
rect 370 184 373 186
rect 365 182 373 184
rect 375 192 382 194
rect 375 190 378 192
rect 380 190 382 192
rect 375 188 382 190
rect 390 193 397 198
rect 390 191 392 193
rect 394 191 397 193
rect 390 189 397 191
rect 375 182 380 188
rect 304 176 307 178
rect 309 176 311 178
rect 304 174 311 176
rect 392 174 397 189
rect 399 185 407 202
rect 399 183 402 185
rect 404 183 407 185
rect 399 178 407 183
rect 399 176 402 178
rect 404 176 407 178
rect 399 174 407 176
rect 409 192 417 202
rect 409 190 412 192
rect 414 190 417 192
rect 409 185 417 190
rect 409 183 412 185
rect 414 183 417 185
rect 409 174 417 183
rect 419 185 426 202
rect 442 200 449 202
rect 442 198 444 200
rect 446 198 449 200
rect 442 193 449 198
rect 442 191 444 193
rect 446 191 449 193
rect 442 189 449 191
rect 419 183 422 185
rect 424 183 426 185
rect 419 178 426 183
rect 419 176 422 178
rect 424 176 426 178
rect 419 174 426 176
rect 444 174 449 189
rect 451 185 459 202
rect 451 183 454 185
rect 456 183 459 185
rect 451 178 459 183
rect 451 176 454 178
rect 456 176 459 178
rect 451 174 459 176
rect 461 192 469 202
rect 461 190 464 192
rect 466 190 469 192
rect 461 185 469 190
rect 461 183 464 185
rect 466 183 469 185
rect 461 174 469 183
rect 471 185 478 202
rect 484 200 491 202
rect 484 198 486 200
rect 488 198 491 200
rect 484 193 491 198
rect 484 191 486 193
rect 488 191 491 193
rect 484 189 491 191
rect 471 183 474 185
rect 476 183 478 185
rect 471 178 478 183
rect 471 176 474 178
rect 476 176 478 178
rect 471 174 478 176
rect 486 174 491 189
rect 493 185 501 202
rect 493 183 496 185
rect 498 183 501 185
rect 493 178 501 183
rect 493 176 496 178
rect 498 176 501 178
rect 493 174 501 176
rect 503 192 511 202
rect 503 190 506 192
rect 508 190 511 192
rect 503 185 511 190
rect 503 183 506 185
rect 508 183 511 185
rect 503 174 511 183
rect 513 185 520 202
rect 528 200 535 202
rect 528 198 530 200
rect 532 198 535 200
rect 528 193 535 198
rect 528 191 530 193
rect 532 191 535 193
rect 528 189 535 191
rect 513 183 516 185
rect 518 183 520 185
rect 513 178 520 183
rect 513 176 516 178
rect 518 176 520 178
rect 513 174 520 176
rect 530 174 535 189
rect 537 185 545 202
rect 537 183 540 185
rect 542 183 545 185
rect 537 178 545 183
rect 537 176 540 178
rect 542 176 545 178
rect 537 174 545 176
rect 547 192 555 202
rect 547 190 550 192
rect 552 190 555 192
rect 547 185 555 190
rect 547 183 550 185
rect 552 183 555 185
rect 547 174 555 183
rect 557 185 564 202
rect 557 183 560 185
rect 562 183 564 185
rect 557 178 564 183
rect 557 176 560 178
rect 562 176 564 178
rect 557 174 564 176
rect 9 150 14 162
rect 7 148 14 150
rect 7 146 9 148
rect 11 146 14 148
rect 7 141 14 146
rect 7 139 9 141
rect 11 139 14 141
rect 7 137 14 139
rect 16 160 25 162
rect 16 158 20 160
rect 22 158 25 160
rect 48 160 62 162
rect 48 159 55 160
rect 16 150 25 158
rect 32 150 37 159
rect 16 137 27 150
rect 29 141 37 150
rect 29 139 32 141
rect 34 139 37 141
rect 29 137 37 139
rect 32 134 37 137
rect 39 134 44 159
rect 46 158 55 159
rect 57 158 62 160
rect 46 153 62 158
rect 46 151 55 153
rect 57 151 62 153
rect 46 134 62 151
rect 64 152 72 162
rect 64 150 67 152
rect 69 150 72 152
rect 64 145 72 150
rect 64 143 67 145
rect 69 143 72 145
rect 64 134 72 143
rect 74 160 82 162
rect 74 158 77 160
rect 79 158 82 160
rect 74 153 82 158
rect 74 151 77 153
rect 79 151 82 153
rect 74 134 82 151
rect 84 147 89 162
rect 105 150 110 162
rect 103 148 110 150
rect 84 145 91 147
rect 84 143 87 145
rect 89 143 91 145
rect 84 138 91 143
rect 84 136 87 138
rect 89 136 91 138
rect 103 146 105 148
rect 107 146 110 148
rect 103 141 110 146
rect 103 139 105 141
rect 107 139 110 141
rect 103 137 110 139
rect 112 160 121 162
rect 112 158 116 160
rect 118 158 121 160
rect 210 163 217 165
rect 210 162 213 163
rect 144 160 158 162
rect 144 159 151 160
rect 112 150 121 158
rect 128 150 133 159
rect 112 137 123 150
rect 125 141 133 150
rect 125 139 128 141
rect 130 139 133 141
rect 125 137 133 139
rect 84 134 91 136
rect 128 134 133 137
rect 135 134 140 159
rect 142 158 151 159
rect 153 158 158 160
rect 142 153 158 158
rect 142 151 151 153
rect 153 151 158 153
rect 142 134 158 151
rect 160 152 168 162
rect 160 150 163 152
rect 165 150 168 152
rect 160 145 168 150
rect 160 143 163 145
rect 165 143 168 145
rect 160 134 168 143
rect 170 160 178 162
rect 170 158 173 160
rect 175 158 178 160
rect 170 153 178 158
rect 170 151 173 153
rect 175 151 178 153
rect 170 134 178 151
rect 180 147 185 162
rect 194 156 199 162
rect 192 154 199 156
rect 192 152 194 154
rect 196 152 199 154
rect 192 150 199 152
rect 180 145 187 147
rect 180 143 183 145
rect 185 143 187 145
rect 180 138 187 143
rect 180 136 183 138
rect 185 136 187 138
rect 180 134 187 136
rect 194 134 199 150
rect 201 134 206 162
rect 208 161 213 162
rect 215 162 217 163
rect 215 161 219 162
rect 208 134 219 161
rect 221 156 226 162
rect 221 154 228 156
rect 221 152 224 154
rect 226 152 228 154
rect 221 147 228 152
rect 249 150 254 162
rect 221 145 224 147
rect 226 145 228 147
rect 221 143 228 145
rect 247 148 254 150
rect 247 146 249 148
rect 251 146 254 148
rect 221 134 226 143
rect 247 141 254 146
rect 247 139 249 141
rect 251 139 254 141
rect 247 137 254 139
rect 256 160 265 162
rect 256 158 260 160
rect 262 158 265 160
rect 288 160 302 162
rect 288 159 295 160
rect 256 150 265 158
rect 272 150 277 159
rect 256 137 267 150
rect 269 141 277 150
rect 269 139 272 141
rect 274 139 277 141
rect 269 137 277 139
rect 272 134 277 137
rect 279 134 284 159
rect 286 158 295 159
rect 297 158 302 160
rect 286 153 302 158
rect 286 151 295 153
rect 297 151 302 153
rect 286 134 302 151
rect 304 152 312 162
rect 304 150 307 152
rect 309 150 312 152
rect 304 145 312 150
rect 304 143 307 145
rect 309 143 312 145
rect 304 134 312 143
rect 314 160 322 162
rect 314 158 317 160
rect 319 158 322 160
rect 314 153 322 158
rect 314 151 317 153
rect 319 151 322 153
rect 314 134 322 151
rect 324 147 329 162
rect 345 150 350 162
rect 343 148 350 150
rect 324 145 331 147
rect 324 143 327 145
rect 329 143 331 145
rect 324 138 331 143
rect 324 136 327 138
rect 329 136 331 138
rect 343 146 345 148
rect 347 146 350 148
rect 343 141 350 146
rect 343 139 345 141
rect 347 139 350 141
rect 343 137 350 139
rect 352 160 361 162
rect 352 158 356 160
rect 358 158 361 160
rect 450 163 457 165
rect 450 162 453 163
rect 384 160 398 162
rect 384 159 391 160
rect 352 150 361 158
rect 368 150 373 159
rect 352 137 363 150
rect 365 141 373 150
rect 365 139 368 141
rect 370 139 373 141
rect 365 137 373 139
rect 324 134 331 136
rect 368 134 373 137
rect 375 134 380 159
rect 382 158 391 159
rect 393 158 398 160
rect 382 153 398 158
rect 382 151 391 153
rect 393 151 398 153
rect 382 134 398 151
rect 400 152 408 162
rect 400 150 403 152
rect 405 150 408 152
rect 400 145 408 150
rect 400 143 403 145
rect 405 143 408 145
rect 400 134 408 143
rect 410 160 418 162
rect 410 158 413 160
rect 415 158 418 160
rect 410 153 418 158
rect 410 151 413 153
rect 415 151 418 153
rect 410 134 418 151
rect 420 147 425 162
rect 434 156 439 162
rect 432 154 439 156
rect 432 152 434 154
rect 436 152 439 154
rect 432 150 439 152
rect 420 145 427 147
rect 420 143 423 145
rect 425 143 427 145
rect 420 138 427 143
rect 420 136 423 138
rect 425 136 427 138
rect 420 134 427 136
rect 434 134 439 150
rect 441 134 446 162
rect 448 161 453 162
rect 455 162 457 163
rect 455 161 459 162
rect 448 134 459 161
rect 461 156 466 162
rect 461 154 468 156
rect 461 152 464 154
rect 466 152 468 154
rect 461 147 468 152
rect 514 152 521 154
rect 514 150 516 152
rect 518 150 521 152
rect 461 145 464 147
rect 466 145 468 147
rect 461 143 468 145
rect 514 148 521 150
rect 461 134 466 143
rect 515 142 521 148
rect 523 142 528 154
rect 530 146 538 154
rect 530 144 533 146
rect 535 144 538 146
rect 530 142 538 144
rect 540 142 545 154
rect 547 152 555 154
rect 547 150 550 152
rect 552 150 555 152
rect 547 142 555 150
rect 557 148 562 154
rect 557 146 564 148
rect 557 144 560 146
rect 562 144 564 146
rect 557 142 564 144
rect 515 140 519 142
rect 504 138 511 140
rect 504 136 506 138
rect 508 136 511 138
rect 504 134 511 136
rect 513 134 519 140
rect 9 49 14 58
rect 7 47 14 49
rect 7 45 9 47
rect 11 45 14 47
rect 7 40 14 45
rect 7 38 9 40
rect 11 38 14 40
rect 7 36 14 38
rect 9 30 14 36
rect 16 31 27 58
rect 16 30 20 31
rect 18 29 20 30
rect 22 30 27 31
rect 29 30 34 58
rect 36 42 41 58
rect 48 56 55 58
rect 48 54 50 56
rect 52 54 55 56
rect 48 49 55 54
rect 48 47 50 49
rect 52 47 55 49
rect 48 45 55 47
rect 36 40 43 42
rect 36 38 39 40
rect 41 38 43 40
rect 36 36 43 38
rect 36 30 41 36
rect 50 30 55 45
rect 57 41 65 58
rect 57 39 60 41
rect 62 39 65 41
rect 57 34 65 39
rect 57 32 60 34
rect 62 32 65 34
rect 57 30 65 32
rect 67 49 75 58
rect 67 47 70 49
rect 72 47 75 49
rect 67 42 75 47
rect 67 40 70 42
rect 72 40 75 42
rect 67 30 75 40
rect 77 41 93 58
rect 77 39 82 41
rect 84 39 93 41
rect 77 34 93 39
rect 77 32 82 34
rect 84 33 93 34
rect 95 33 100 58
rect 102 55 107 58
rect 144 56 151 58
rect 102 53 110 55
rect 102 51 105 53
rect 107 51 110 53
rect 102 42 110 51
rect 112 42 123 55
rect 102 33 107 42
rect 114 34 123 42
rect 84 32 91 33
rect 77 30 91 32
rect 22 29 25 30
rect 18 27 25 29
rect 114 32 117 34
rect 119 32 123 34
rect 114 30 123 32
rect 125 53 132 55
rect 125 51 128 53
rect 130 51 132 53
rect 125 46 132 51
rect 125 44 128 46
rect 130 44 132 46
rect 144 54 146 56
rect 148 54 151 56
rect 144 49 151 54
rect 144 47 146 49
rect 148 47 151 49
rect 144 45 151 47
rect 125 42 132 44
rect 125 30 130 42
rect 146 30 151 45
rect 153 41 161 58
rect 153 39 156 41
rect 158 39 161 41
rect 153 34 161 39
rect 153 32 156 34
rect 158 32 161 34
rect 153 30 161 32
rect 163 49 171 58
rect 163 47 166 49
rect 168 47 171 49
rect 163 42 171 47
rect 163 40 166 42
rect 168 40 171 42
rect 163 30 171 40
rect 173 41 189 58
rect 173 39 178 41
rect 180 39 189 41
rect 173 34 189 39
rect 173 32 178 34
rect 180 33 189 34
rect 191 33 196 58
rect 198 55 203 58
rect 198 53 206 55
rect 198 51 201 53
rect 203 51 206 53
rect 198 42 206 51
rect 208 42 219 55
rect 198 33 203 42
rect 210 34 219 42
rect 180 32 187 33
rect 173 30 187 32
rect 210 32 213 34
rect 215 32 219 34
rect 210 30 219 32
rect 221 53 228 55
rect 221 51 224 53
rect 226 51 228 53
rect 221 46 228 51
rect 248 49 253 58
rect 221 44 224 46
rect 226 44 228 46
rect 221 42 228 44
rect 246 47 253 49
rect 246 45 248 47
rect 250 45 253 47
rect 221 30 226 42
rect 246 40 253 45
rect 246 38 248 40
rect 250 38 253 40
rect 246 36 253 38
rect 248 30 253 36
rect 255 31 266 58
rect 255 30 259 31
rect 257 29 259 30
rect 261 30 266 31
rect 268 30 273 58
rect 275 42 280 58
rect 287 56 294 58
rect 287 54 289 56
rect 291 54 294 56
rect 287 49 294 54
rect 287 47 289 49
rect 291 47 294 49
rect 287 45 294 47
rect 275 40 282 42
rect 275 38 278 40
rect 280 38 282 40
rect 275 36 282 38
rect 275 30 280 36
rect 289 30 294 45
rect 296 41 304 58
rect 296 39 299 41
rect 301 39 304 41
rect 296 34 304 39
rect 296 32 299 34
rect 301 32 304 34
rect 296 30 304 32
rect 306 49 314 58
rect 306 47 309 49
rect 311 47 314 49
rect 306 42 314 47
rect 306 40 309 42
rect 311 40 314 42
rect 306 30 314 40
rect 316 41 332 58
rect 316 39 321 41
rect 323 39 332 41
rect 316 34 332 39
rect 316 32 321 34
rect 323 33 332 34
rect 334 33 339 58
rect 341 55 346 58
rect 383 56 390 58
rect 341 53 349 55
rect 341 51 344 53
rect 346 51 349 53
rect 341 42 349 51
rect 351 42 362 55
rect 341 33 346 42
rect 353 34 362 42
rect 323 32 330 33
rect 316 30 330 32
rect 261 29 264 30
rect 257 27 264 29
rect 353 32 356 34
rect 358 32 362 34
rect 353 30 362 32
rect 364 53 371 55
rect 364 51 367 53
rect 369 51 371 53
rect 364 46 371 51
rect 364 44 367 46
rect 369 44 371 46
rect 383 54 385 56
rect 387 54 390 56
rect 383 49 390 54
rect 383 47 385 49
rect 387 47 390 49
rect 383 45 390 47
rect 364 42 371 44
rect 364 30 369 42
rect 385 30 390 45
rect 392 41 400 58
rect 392 39 395 41
rect 397 39 400 41
rect 392 34 400 39
rect 392 32 395 34
rect 397 32 400 34
rect 392 30 400 32
rect 402 49 410 58
rect 402 47 405 49
rect 407 47 410 49
rect 402 42 410 47
rect 402 40 405 42
rect 407 40 410 42
rect 402 30 410 40
rect 412 41 428 58
rect 412 39 417 41
rect 419 39 428 41
rect 412 34 428 39
rect 412 32 417 34
rect 419 33 428 34
rect 430 33 435 58
rect 437 55 442 58
rect 504 56 511 58
rect 437 53 445 55
rect 437 51 440 53
rect 442 51 445 53
rect 437 42 445 51
rect 447 42 458 55
rect 437 33 442 42
rect 449 34 458 42
rect 419 32 426 33
rect 412 30 426 32
rect 449 32 452 34
rect 454 32 458 34
rect 449 30 458 32
rect 460 53 467 55
rect 460 51 463 53
rect 465 51 467 53
rect 504 54 506 56
rect 508 54 511 56
rect 504 52 511 54
rect 513 52 519 58
rect 460 46 467 51
rect 460 44 463 46
rect 465 44 467 46
rect 460 42 467 44
rect 515 50 519 52
rect 515 44 521 50
rect 514 42 521 44
rect 460 30 465 42
rect 514 40 516 42
rect 518 40 521 42
rect 514 38 521 40
rect 523 38 528 50
rect 530 48 538 50
rect 530 46 533 48
rect 535 46 538 48
rect 530 38 538 46
rect 540 38 545 50
rect 547 42 555 50
rect 547 40 550 42
rect 552 40 555 42
rect 547 38 555 40
rect 557 48 564 50
rect 557 46 560 48
rect 562 46 564 48
rect 557 44 564 46
rect 557 38 562 44
rect 9 6 14 18
rect 7 4 14 6
rect 7 2 9 4
rect 11 2 14 4
rect 7 -3 14 2
rect 7 -5 9 -3
rect 11 -5 14 -3
rect 7 -7 14 -5
rect 16 16 25 18
rect 16 14 20 16
rect 22 14 25 16
rect 48 16 62 18
rect 48 15 55 16
rect 16 6 25 14
rect 32 6 37 15
rect 16 -7 27 6
rect 29 -3 37 6
rect 29 -5 32 -3
rect 34 -5 37 -3
rect 29 -7 37 -5
rect 32 -10 37 -7
rect 39 -10 44 15
rect 46 14 55 15
rect 57 14 62 16
rect 46 9 62 14
rect 46 7 55 9
rect 57 7 62 9
rect 46 -10 62 7
rect 64 8 72 18
rect 64 6 67 8
rect 69 6 72 8
rect 64 1 72 6
rect 64 -1 67 1
rect 69 -1 72 1
rect 64 -10 72 -1
rect 74 16 82 18
rect 74 14 77 16
rect 79 14 82 16
rect 74 9 82 14
rect 74 7 77 9
rect 79 7 82 9
rect 74 -10 82 7
rect 84 3 89 18
rect 105 6 110 18
rect 103 4 110 6
rect 84 1 91 3
rect 84 -1 87 1
rect 89 -1 91 1
rect 84 -6 91 -1
rect 84 -8 87 -6
rect 89 -8 91 -6
rect 103 2 105 4
rect 107 2 110 4
rect 103 -3 110 2
rect 103 -5 105 -3
rect 107 -5 110 -3
rect 103 -7 110 -5
rect 112 16 121 18
rect 112 14 116 16
rect 118 14 121 16
rect 210 19 217 21
rect 210 18 213 19
rect 144 16 158 18
rect 144 15 151 16
rect 112 6 121 14
rect 128 6 133 15
rect 112 -7 123 6
rect 125 -3 133 6
rect 125 -5 128 -3
rect 130 -5 133 -3
rect 125 -7 133 -5
rect 84 -10 91 -8
rect 128 -10 133 -7
rect 135 -10 140 15
rect 142 14 151 15
rect 153 14 158 16
rect 142 9 158 14
rect 142 7 151 9
rect 153 7 158 9
rect 142 -10 158 7
rect 160 8 168 18
rect 160 6 163 8
rect 165 6 168 8
rect 160 1 168 6
rect 160 -1 163 1
rect 165 -1 168 1
rect 160 -10 168 -1
rect 170 16 178 18
rect 170 14 173 16
rect 175 14 178 16
rect 170 9 178 14
rect 170 7 173 9
rect 175 7 178 9
rect 170 -10 178 7
rect 180 3 185 18
rect 194 12 199 18
rect 192 10 199 12
rect 192 8 194 10
rect 196 8 199 10
rect 192 6 199 8
rect 180 1 187 3
rect 180 -1 183 1
rect 185 -1 187 1
rect 180 -6 187 -1
rect 180 -8 183 -6
rect 185 -8 187 -6
rect 180 -10 187 -8
rect 194 -10 199 6
rect 201 -10 206 18
rect 208 17 213 18
rect 215 18 217 19
rect 215 17 219 18
rect 208 -10 219 17
rect 221 12 226 18
rect 221 10 228 12
rect 221 8 224 10
rect 226 8 228 10
rect 221 3 228 8
rect 249 6 254 18
rect 221 1 224 3
rect 226 1 228 3
rect 221 -1 228 1
rect 247 4 254 6
rect 247 2 249 4
rect 251 2 254 4
rect 221 -10 226 -1
rect 247 -3 254 2
rect 247 -5 249 -3
rect 251 -5 254 -3
rect 247 -7 254 -5
rect 256 16 265 18
rect 256 14 260 16
rect 262 14 265 16
rect 288 16 302 18
rect 288 15 295 16
rect 256 6 265 14
rect 272 6 277 15
rect 256 -7 267 6
rect 269 -3 277 6
rect 269 -5 272 -3
rect 274 -5 277 -3
rect 269 -7 277 -5
rect 272 -10 277 -7
rect 279 -10 284 15
rect 286 14 295 15
rect 297 14 302 16
rect 286 9 302 14
rect 286 7 295 9
rect 297 7 302 9
rect 286 -10 302 7
rect 304 8 312 18
rect 304 6 307 8
rect 309 6 312 8
rect 304 1 312 6
rect 304 -1 307 1
rect 309 -1 312 1
rect 304 -10 312 -1
rect 314 16 322 18
rect 314 14 317 16
rect 319 14 322 16
rect 314 9 322 14
rect 314 7 317 9
rect 319 7 322 9
rect 314 -10 322 7
rect 324 3 329 18
rect 345 6 350 18
rect 343 4 350 6
rect 324 1 331 3
rect 324 -1 327 1
rect 329 -1 331 1
rect 324 -6 331 -1
rect 324 -8 327 -6
rect 329 -8 331 -6
rect 343 2 345 4
rect 347 2 350 4
rect 343 -3 350 2
rect 343 -5 345 -3
rect 347 -5 350 -3
rect 343 -7 350 -5
rect 352 16 361 18
rect 352 14 356 16
rect 358 14 361 16
rect 450 19 457 21
rect 450 18 453 19
rect 384 16 398 18
rect 384 15 391 16
rect 352 6 361 14
rect 368 6 373 15
rect 352 -7 363 6
rect 365 -3 373 6
rect 365 -5 368 -3
rect 370 -5 373 -3
rect 365 -7 373 -5
rect 324 -10 331 -8
rect 368 -10 373 -7
rect 375 -10 380 15
rect 382 14 391 15
rect 393 14 398 16
rect 382 9 398 14
rect 382 7 391 9
rect 393 7 398 9
rect 382 -10 398 7
rect 400 8 408 18
rect 400 6 403 8
rect 405 6 408 8
rect 400 1 408 6
rect 400 -1 403 1
rect 405 -1 408 1
rect 400 -10 408 -1
rect 410 16 418 18
rect 410 14 413 16
rect 415 14 418 16
rect 410 9 418 14
rect 410 7 413 9
rect 415 7 418 9
rect 410 -10 418 7
rect 420 3 425 18
rect 434 12 439 18
rect 432 10 439 12
rect 432 8 434 10
rect 436 8 439 10
rect 432 6 439 8
rect 420 1 427 3
rect 420 -1 423 1
rect 425 -1 427 1
rect 420 -6 427 -1
rect 420 -8 423 -6
rect 425 -8 427 -6
rect 420 -10 427 -8
rect 434 -10 439 6
rect 441 -10 446 18
rect 448 17 453 18
rect 455 18 457 19
rect 455 17 459 18
rect 448 -10 459 17
rect 461 12 466 18
rect 461 10 468 12
rect 461 8 464 10
rect 466 8 468 10
rect 461 3 468 8
rect 514 8 521 10
rect 514 6 516 8
rect 518 6 521 8
rect 461 1 464 3
rect 466 1 468 3
rect 461 -1 468 1
rect 514 4 521 6
rect 461 -10 466 -1
rect 515 -2 521 4
rect 523 -2 528 10
rect 530 2 538 10
rect 530 0 533 2
rect 535 0 538 2
rect 530 -2 538 0
rect 540 -2 545 10
rect 547 8 555 10
rect 547 6 550 8
rect 552 6 555 8
rect 547 -2 555 6
rect 557 4 562 10
rect 557 2 564 4
rect 557 0 560 2
rect 562 0 564 2
rect 557 -2 564 0
rect 515 -4 519 -2
rect 504 -6 511 -4
rect 504 -8 506 -6
rect 508 -8 511 -6
rect 504 -10 511 -8
rect 513 -10 519 -4
rect 9 -95 14 -86
rect 7 -97 14 -95
rect 7 -99 9 -97
rect 11 -99 14 -97
rect 7 -104 14 -99
rect 7 -106 9 -104
rect 11 -106 14 -104
rect 7 -108 14 -106
rect 9 -114 14 -108
rect 16 -113 27 -86
rect 16 -114 20 -113
rect 18 -115 20 -114
rect 22 -114 27 -113
rect 29 -114 34 -86
rect 36 -102 41 -86
rect 48 -88 55 -86
rect 48 -90 50 -88
rect 52 -90 55 -88
rect 48 -95 55 -90
rect 48 -97 50 -95
rect 52 -97 55 -95
rect 48 -99 55 -97
rect 36 -104 43 -102
rect 36 -106 39 -104
rect 41 -106 43 -104
rect 36 -108 43 -106
rect 36 -114 41 -108
rect 50 -114 55 -99
rect 57 -103 65 -86
rect 57 -105 60 -103
rect 62 -105 65 -103
rect 57 -110 65 -105
rect 57 -112 60 -110
rect 62 -112 65 -110
rect 57 -114 65 -112
rect 67 -95 75 -86
rect 67 -97 70 -95
rect 72 -97 75 -95
rect 67 -102 75 -97
rect 67 -104 70 -102
rect 72 -104 75 -102
rect 67 -114 75 -104
rect 77 -103 93 -86
rect 77 -105 82 -103
rect 84 -105 93 -103
rect 77 -110 93 -105
rect 77 -112 82 -110
rect 84 -111 93 -110
rect 95 -111 100 -86
rect 102 -89 107 -86
rect 144 -88 151 -86
rect 102 -91 110 -89
rect 102 -93 105 -91
rect 107 -93 110 -91
rect 102 -102 110 -93
rect 112 -102 123 -89
rect 102 -111 107 -102
rect 114 -110 123 -102
rect 84 -112 91 -111
rect 77 -114 91 -112
rect 22 -115 25 -114
rect 18 -117 25 -115
rect 114 -112 117 -110
rect 119 -112 123 -110
rect 114 -114 123 -112
rect 125 -91 132 -89
rect 125 -93 128 -91
rect 130 -93 132 -91
rect 125 -98 132 -93
rect 125 -100 128 -98
rect 130 -100 132 -98
rect 144 -90 146 -88
rect 148 -90 151 -88
rect 144 -95 151 -90
rect 144 -97 146 -95
rect 148 -97 151 -95
rect 144 -99 151 -97
rect 125 -102 132 -100
rect 125 -114 130 -102
rect 146 -114 151 -99
rect 153 -103 161 -86
rect 153 -105 156 -103
rect 158 -105 161 -103
rect 153 -110 161 -105
rect 153 -112 156 -110
rect 158 -112 161 -110
rect 153 -114 161 -112
rect 163 -95 171 -86
rect 163 -97 166 -95
rect 168 -97 171 -95
rect 163 -102 171 -97
rect 163 -104 166 -102
rect 168 -104 171 -102
rect 163 -114 171 -104
rect 173 -103 189 -86
rect 173 -105 178 -103
rect 180 -105 189 -103
rect 173 -110 189 -105
rect 173 -112 178 -110
rect 180 -111 189 -110
rect 191 -111 196 -86
rect 198 -89 203 -86
rect 198 -91 206 -89
rect 198 -93 201 -91
rect 203 -93 206 -91
rect 198 -102 206 -93
rect 208 -102 219 -89
rect 198 -111 203 -102
rect 210 -110 219 -102
rect 180 -112 187 -111
rect 173 -114 187 -112
rect 210 -112 213 -110
rect 215 -112 219 -110
rect 210 -114 219 -112
rect 221 -91 228 -89
rect 221 -93 224 -91
rect 226 -93 228 -91
rect 221 -98 228 -93
rect 248 -95 253 -86
rect 221 -100 224 -98
rect 226 -100 228 -98
rect 221 -102 228 -100
rect 246 -97 253 -95
rect 246 -99 248 -97
rect 250 -99 253 -97
rect 221 -114 226 -102
rect 246 -104 253 -99
rect 246 -106 248 -104
rect 250 -106 253 -104
rect 246 -108 253 -106
rect 248 -114 253 -108
rect 255 -113 266 -86
rect 255 -114 259 -113
rect 257 -115 259 -114
rect 261 -114 266 -113
rect 268 -114 273 -86
rect 275 -102 280 -86
rect 287 -88 294 -86
rect 287 -90 289 -88
rect 291 -90 294 -88
rect 287 -95 294 -90
rect 287 -97 289 -95
rect 291 -97 294 -95
rect 287 -99 294 -97
rect 275 -104 282 -102
rect 275 -106 278 -104
rect 280 -106 282 -104
rect 275 -108 282 -106
rect 275 -114 280 -108
rect 289 -114 294 -99
rect 296 -103 304 -86
rect 296 -105 299 -103
rect 301 -105 304 -103
rect 296 -110 304 -105
rect 296 -112 299 -110
rect 301 -112 304 -110
rect 296 -114 304 -112
rect 306 -95 314 -86
rect 306 -97 309 -95
rect 311 -97 314 -95
rect 306 -102 314 -97
rect 306 -104 309 -102
rect 311 -104 314 -102
rect 306 -114 314 -104
rect 316 -103 332 -86
rect 316 -105 321 -103
rect 323 -105 332 -103
rect 316 -110 332 -105
rect 316 -112 321 -110
rect 323 -111 332 -110
rect 334 -111 339 -86
rect 341 -89 346 -86
rect 383 -88 390 -86
rect 341 -91 349 -89
rect 341 -93 344 -91
rect 346 -93 349 -91
rect 341 -102 349 -93
rect 351 -102 362 -89
rect 341 -111 346 -102
rect 353 -110 362 -102
rect 323 -112 330 -111
rect 316 -114 330 -112
rect 261 -115 264 -114
rect 257 -117 264 -115
rect 353 -112 356 -110
rect 358 -112 362 -110
rect 353 -114 362 -112
rect 364 -91 371 -89
rect 364 -93 367 -91
rect 369 -93 371 -91
rect 364 -98 371 -93
rect 364 -100 367 -98
rect 369 -100 371 -98
rect 383 -90 385 -88
rect 387 -90 390 -88
rect 383 -95 390 -90
rect 383 -97 385 -95
rect 387 -97 390 -95
rect 383 -99 390 -97
rect 364 -102 371 -100
rect 364 -114 369 -102
rect 385 -114 390 -99
rect 392 -103 400 -86
rect 392 -105 395 -103
rect 397 -105 400 -103
rect 392 -110 400 -105
rect 392 -112 395 -110
rect 397 -112 400 -110
rect 392 -114 400 -112
rect 402 -95 410 -86
rect 402 -97 405 -95
rect 407 -97 410 -95
rect 402 -102 410 -97
rect 402 -104 405 -102
rect 407 -104 410 -102
rect 402 -114 410 -104
rect 412 -103 428 -86
rect 412 -105 417 -103
rect 419 -105 428 -103
rect 412 -110 428 -105
rect 412 -112 417 -110
rect 419 -111 428 -110
rect 430 -111 435 -86
rect 437 -89 442 -86
rect 504 -88 511 -86
rect 437 -91 445 -89
rect 437 -93 440 -91
rect 442 -93 445 -91
rect 437 -102 445 -93
rect 447 -102 458 -89
rect 437 -111 442 -102
rect 449 -110 458 -102
rect 419 -112 426 -111
rect 412 -114 426 -112
rect 449 -112 452 -110
rect 454 -112 458 -110
rect 449 -114 458 -112
rect 460 -91 467 -89
rect 460 -93 463 -91
rect 465 -93 467 -91
rect 504 -90 506 -88
rect 508 -90 511 -88
rect 504 -92 511 -90
rect 513 -92 519 -86
rect 460 -98 467 -93
rect 460 -100 463 -98
rect 465 -100 467 -98
rect 460 -102 467 -100
rect 515 -94 519 -92
rect 515 -100 521 -94
rect 514 -102 521 -100
rect 460 -114 465 -102
rect 514 -104 516 -102
rect 518 -104 521 -102
rect 514 -106 521 -104
rect 523 -106 528 -94
rect 530 -96 538 -94
rect 530 -98 533 -96
rect 535 -98 538 -96
rect 530 -106 538 -98
rect 540 -106 545 -94
rect 547 -102 555 -94
rect 547 -104 550 -102
rect 552 -104 555 -102
rect 547 -106 555 -104
rect 557 -96 564 -94
rect 557 -98 560 -96
rect 562 -98 564 -96
rect 557 -100 564 -98
rect 557 -106 562 -100
<< alu1 >>
rect 3 235 568 240
rect 3 233 86 235
rect 88 233 109 235
rect 111 233 119 235
rect 121 233 127 235
rect 129 233 286 235
rect 288 233 568 235
rect 3 232 568 233
rect 24 225 28 227
rect 26 223 28 225
rect 24 218 28 223
rect 26 216 28 218
rect 8 209 20 211
rect 8 207 16 209
rect 18 207 20 209
rect 8 205 20 207
rect 24 205 28 216
rect 57 225 61 227
rect 59 223 61 225
rect 57 218 61 223
rect 59 216 61 218
rect 8 189 12 205
rect 24 203 25 205
rect 27 203 28 205
rect 24 199 28 203
rect 26 197 28 199
rect 24 195 28 197
rect 16 192 28 195
rect 16 190 24 192
rect 26 190 28 192
rect 16 189 28 190
rect 41 209 53 211
rect 41 207 49 209
rect 51 207 53 209
rect 41 205 53 207
rect 41 189 45 205
rect 57 199 61 216
rect 87 218 92 227
rect 96 225 121 226
rect 96 223 98 225
rect 100 223 121 225
rect 96 222 118 223
rect 117 221 118 222
rect 120 221 121 223
rect 87 217 109 218
rect 87 215 88 217
rect 90 216 109 217
rect 90 215 101 216
rect 87 214 101 215
rect 103 214 109 216
rect 117 214 121 221
rect 146 225 150 227
rect 146 223 148 225
rect 146 218 150 223
rect 146 216 148 218
rect 59 197 61 199
rect 88 209 101 210
rect 88 207 89 209
rect 91 207 101 209
rect 88 206 101 207
rect 117 210 132 214
rect 88 203 92 206
rect 88 201 89 203
rect 91 201 92 203
rect 88 197 92 201
rect 96 198 112 202
rect 120 203 124 205
rect 120 201 121 203
rect 123 201 124 203
rect 57 195 61 197
rect 49 193 61 195
rect 49 192 67 193
rect 49 190 57 192
rect 59 190 64 192
rect 66 190 67 192
rect 49 189 67 190
rect 96 184 100 198
rect 120 194 124 201
rect 111 193 124 194
rect 111 191 117 193
rect 119 191 124 193
rect 111 190 124 191
rect 128 186 132 210
rect 146 199 150 216
rect 194 225 198 227
rect 196 223 198 225
rect 194 218 198 223
rect 196 216 198 218
rect 154 209 166 211
rect 154 207 156 209
rect 158 207 166 209
rect 154 205 166 207
rect 146 197 148 199
rect 146 195 150 197
rect 146 193 158 195
rect 142 192 158 193
rect 142 190 143 192
rect 145 190 148 192
rect 150 190 158 192
rect 142 189 158 190
rect 162 189 166 205
rect 178 209 190 211
rect 178 207 186 209
rect 188 207 190 209
rect 178 205 190 207
rect 178 189 182 205
rect 194 199 198 216
rect 196 197 198 199
rect 266 226 272 227
rect 266 224 268 226
rect 270 224 272 226
rect 266 223 272 224
rect 220 213 232 219
rect 226 209 232 213
rect 226 207 227 209
rect 229 207 232 209
rect 226 205 232 207
rect 243 207 258 210
rect 243 205 254 207
rect 256 205 258 207
rect 243 204 258 205
rect 243 201 249 204
rect 243 199 246 201
rect 248 199 249 201
rect 243 198 249 199
rect 268 211 272 223
rect 295 218 311 219
rect 295 216 297 218
rect 299 216 311 218
rect 295 215 311 216
rect 268 209 296 211
rect 268 207 293 209
rect 295 207 296 209
rect 268 205 296 207
rect 194 195 200 197
rect 186 193 197 195
rect 199 193 200 195
rect 268 194 272 205
rect 290 198 296 205
rect 307 201 311 215
rect 307 199 308 201
rect 310 199 311 201
rect 307 194 311 199
rect 376 226 382 227
rect 376 224 378 226
rect 380 224 382 226
rect 376 223 382 224
rect 330 213 342 219
rect 336 209 342 213
rect 336 207 337 209
rect 339 207 342 209
rect 336 205 342 207
rect 353 207 368 210
rect 353 205 364 207
rect 366 205 368 207
rect 353 204 368 205
rect 353 201 359 204
rect 353 199 354 201
rect 356 199 359 201
rect 353 198 359 199
rect 378 194 382 223
rect 186 192 200 193
rect 186 190 194 192
rect 196 190 198 192
rect 186 189 198 190
rect 212 191 225 194
rect 212 189 214 191
rect 216 190 225 191
rect 259 192 272 194
rect 259 190 268 192
rect 270 190 272 192
rect 290 192 311 194
rect 290 190 297 192
rect 299 190 311 192
rect 322 191 335 194
rect 216 189 217 190
rect 266 189 272 190
rect 96 182 97 184
rect 99 182 100 184
rect 96 181 100 182
rect 117 185 132 186
rect 117 183 119 185
rect 121 184 132 185
rect 121 183 129 184
rect 117 182 129 183
rect 131 182 132 184
rect 117 181 132 182
rect 212 184 217 189
rect 212 182 213 184
rect 215 182 217 184
rect 212 181 217 182
rect 322 189 324 191
rect 326 190 335 191
rect 369 192 382 194
rect 369 190 378 192
rect 380 190 382 192
rect 326 189 327 190
rect 376 189 382 190
rect 411 225 418 227
rect 411 223 412 225
rect 414 223 418 225
rect 411 221 418 223
rect 397 209 402 211
rect 397 207 398 209
rect 400 207 402 209
rect 397 205 402 207
rect 414 211 418 221
rect 463 225 470 227
rect 463 223 464 225
rect 466 223 470 225
rect 463 221 470 223
rect 414 207 426 211
rect 398 202 402 205
rect 398 198 411 202
rect 422 194 426 207
rect 411 193 426 194
rect 411 192 423 193
rect 411 190 412 192
rect 414 191 423 192
rect 425 191 426 193
rect 414 190 426 191
rect 449 209 454 211
rect 449 207 450 209
rect 452 207 454 209
rect 449 205 454 207
rect 466 211 470 221
rect 505 225 512 227
rect 505 223 506 225
rect 508 223 512 225
rect 505 221 512 223
rect 466 207 478 211
rect 450 202 454 205
rect 450 198 463 202
rect 474 194 478 207
rect 322 184 327 189
rect 322 182 323 184
rect 325 182 327 184
rect 322 181 327 182
rect 411 185 415 190
rect 463 193 478 194
rect 463 192 475 193
rect 463 190 464 192
rect 466 191 475 192
rect 477 191 478 193
rect 466 190 478 191
rect 491 209 496 211
rect 491 207 492 209
rect 494 207 496 209
rect 491 205 496 207
rect 508 211 512 221
rect 549 225 556 227
rect 549 223 550 225
rect 552 223 556 225
rect 549 221 556 223
rect 508 207 520 211
rect 492 202 496 205
rect 492 198 505 202
rect 516 194 520 207
rect 411 183 412 185
rect 414 183 415 185
rect 411 181 415 183
rect 463 185 467 190
rect 505 193 520 194
rect 505 192 517 193
rect 505 190 506 192
rect 508 191 517 192
rect 519 191 520 193
rect 508 190 520 191
rect 535 209 540 211
rect 535 207 536 209
rect 538 207 540 209
rect 535 205 540 207
rect 552 211 556 221
rect 552 207 564 211
rect 536 202 540 205
rect 536 198 549 202
rect 560 194 564 207
rect 463 183 464 185
rect 466 183 467 185
rect 463 181 467 183
rect 505 185 509 190
rect 549 193 564 194
rect 549 192 561 193
rect 549 190 550 192
rect 552 191 561 192
rect 563 191 564 193
rect 552 190 564 191
rect 505 183 506 185
rect 508 183 509 185
rect 505 181 509 183
rect 549 185 553 190
rect 549 183 550 185
rect 552 183 553 185
rect 549 181 553 183
rect 3 175 568 176
rect 3 173 127 175
rect 129 173 215 175
rect 217 173 325 175
rect 327 173 568 175
rect 3 163 568 173
rect 3 161 213 163
rect 215 161 453 163
rect 455 161 507 163
rect 509 161 568 163
rect 3 160 568 161
rect 7 153 20 154
rect 7 151 8 153
rect 10 151 20 153
rect 7 150 20 151
rect 103 150 116 154
rect 7 148 12 150
rect 7 146 9 148
rect 11 146 12 148
rect 103 148 108 150
rect 7 141 12 146
rect 7 139 9 141
rect 11 139 12 141
rect 7 137 12 139
rect 7 115 11 137
rect 38 134 76 138
rect 38 131 43 134
rect 35 129 43 131
rect 35 127 36 129
rect 38 127 43 129
rect 35 125 43 127
rect 53 129 68 130
rect 53 127 55 129
rect 57 127 62 129
rect 64 127 68 129
rect 53 126 68 127
rect 55 122 59 126
rect 86 145 92 147
rect 86 143 87 145
rect 89 143 92 145
rect 86 138 92 143
rect 86 136 87 138
rect 89 136 92 138
rect 86 134 92 136
rect 7 113 12 115
rect 55 120 56 122
rect 58 120 59 122
rect 55 117 59 120
rect 88 115 92 134
rect 103 146 105 148
rect 107 146 108 148
rect 103 141 108 146
rect 103 139 105 141
rect 107 139 108 141
rect 103 137 108 139
rect 103 122 107 137
rect 134 137 172 138
rect 134 135 151 137
rect 153 135 172 137
rect 134 134 172 135
rect 134 131 139 134
rect 131 129 139 131
rect 131 127 132 129
rect 134 127 139 129
rect 131 125 139 127
rect 149 129 164 130
rect 149 127 151 129
rect 153 127 158 129
rect 160 127 164 129
rect 149 126 164 127
rect 103 120 104 122
rect 106 120 107 122
rect 103 115 107 120
rect 88 114 99 115
rect 7 111 9 113
rect 11 111 12 113
rect 7 109 12 111
rect 70 113 99 114
rect 70 111 87 113
rect 89 111 96 113
rect 98 111 99 113
rect 70 110 99 111
rect 103 113 108 115
rect 151 117 155 126
rect 182 145 204 147
rect 182 143 183 145
rect 185 143 204 145
rect 182 141 204 143
rect 216 154 228 155
rect 216 152 224 154
rect 226 152 228 154
rect 216 149 228 152
rect 224 147 228 149
rect 226 145 228 147
rect 182 138 188 141
rect 182 136 183 138
rect 185 136 188 138
rect 182 134 188 136
rect 184 114 188 134
rect 192 129 196 141
rect 192 127 194 129
rect 192 125 196 127
rect 208 138 212 139
rect 208 136 209 138
rect 211 136 212 138
rect 208 131 212 136
rect 200 129 212 131
rect 200 127 207 129
rect 209 127 212 129
rect 200 125 212 127
rect 224 133 228 145
rect 247 150 260 154
rect 343 150 356 154
rect 247 148 252 150
rect 247 146 249 148
rect 251 146 252 148
rect 343 148 348 150
rect 247 141 252 146
rect 247 139 249 141
rect 251 139 252 141
rect 247 137 252 139
rect 224 132 243 133
rect 224 130 240 132
rect 242 130 243 132
rect 224 129 243 130
rect 224 122 228 129
rect 223 120 228 122
rect 223 118 224 120
rect 226 118 228 120
rect 103 111 105 113
rect 107 111 108 113
rect 103 109 108 111
rect 166 113 188 114
rect 166 111 183 113
rect 185 111 188 113
rect 166 110 188 111
rect 223 113 228 118
rect 223 111 224 113
rect 226 111 228 113
rect 223 109 228 111
rect 247 124 251 137
rect 278 134 316 138
rect 247 122 248 124
rect 250 122 251 124
rect 278 132 283 134
rect 278 131 280 132
rect 275 130 280 131
rect 282 130 283 132
rect 275 129 283 130
rect 275 127 276 129
rect 278 127 283 129
rect 275 125 283 127
rect 293 129 308 130
rect 293 127 295 129
rect 297 127 302 129
rect 304 127 308 129
rect 293 126 308 127
rect 247 115 251 122
rect 295 122 299 126
rect 326 145 332 147
rect 326 143 327 145
rect 329 143 332 145
rect 326 138 332 143
rect 326 136 327 138
rect 329 136 332 138
rect 326 134 332 136
rect 247 113 252 115
rect 295 120 296 122
rect 298 120 299 122
rect 295 117 299 120
rect 328 115 332 134
rect 343 146 345 148
rect 347 146 348 148
rect 343 141 348 146
rect 343 139 345 141
rect 347 139 348 141
rect 343 137 348 139
rect 343 122 347 137
rect 374 137 412 138
rect 374 135 376 137
rect 378 135 412 137
rect 374 134 412 135
rect 374 131 379 134
rect 371 129 379 131
rect 371 127 372 129
rect 374 127 379 129
rect 371 125 379 127
rect 389 129 404 130
rect 389 127 391 129
rect 393 127 398 129
rect 400 127 404 129
rect 389 126 404 127
rect 343 120 344 122
rect 346 120 347 122
rect 343 115 347 120
rect 328 114 339 115
rect 247 111 249 113
rect 251 111 252 113
rect 247 109 252 111
rect 310 113 339 114
rect 310 111 327 113
rect 329 111 336 113
rect 338 111 339 113
rect 310 110 339 111
rect 343 113 348 115
rect 391 117 395 126
rect 422 145 444 147
rect 422 143 423 145
rect 425 143 444 145
rect 422 141 444 143
rect 456 154 468 155
rect 456 152 464 154
rect 466 152 468 154
rect 456 149 468 152
rect 464 147 468 149
rect 466 145 468 147
rect 422 138 428 141
rect 422 136 423 138
rect 425 136 428 138
rect 422 134 428 136
rect 424 114 428 134
rect 432 129 436 141
rect 432 127 434 129
rect 432 125 436 127
rect 448 138 452 139
rect 448 136 449 138
rect 451 136 452 138
rect 448 131 452 136
rect 440 129 452 131
rect 440 127 447 129
rect 449 127 452 129
rect 440 125 452 127
rect 464 133 468 145
rect 504 147 509 155
rect 504 145 506 147
rect 508 146 509 147
rect 558 146 564 147
rect 508 145 517 146
rect 504 142 517 145
rect 551 144 560 146
rect 562 144 564 146
rect 551 142 564 144
rect 464 132 484 133
rect 464 130 481 132
rect 483 130 484 132
rect 464 129 484 130
rect 464 122 468 129
rect 463 120 468 122
rect 463 118 464 120
rect 466 118 468 120
rect 343 111 345 113
rect 347 111 348 113
rect 343 109 348 111
rect 406 113 428 114
rect 406 111 423 113
rect 425 111 428 113
rect 406 110 428 111
rect 463 113 468 118
rect 463 111 464 113
rect 466 111 468 113
rect 463 109 468 111
rect 518 129 524 131
rect 518 127 519 129
rect 521 127 524 129
rect 518 123 524 127
rect 512 122 524 123
rect 512 120 514 122
rect 516 120 524 122
rect 512 117 524 120
rect 535 132 541 138
rect 535 131 550 132
rect 535 129 546 131
rect 548 129 550 131
rect 535 126 550 129
rect 560 113 564 142
rect 558 112 564 113
rect 558 110 560 112
rect 562 110 564 112
rect 558 109 564 110
rect 3 103 568 104
rect 3 101 197 103
rect 199 101 437 103
rect 439 101 568 103
rect 3 91 568 101
rect 3 89 36 91
rect 38 89 275 91
rect 277 89 568 91
rect 3 88 568 89
rect 7 81 12 83
rect 7 79 9 81
rect 11 79 12 81
rect 7 74 12 79
rect 47 81 69 82
rect 47 79 50 81
rect 52 79 69 81
rect 47 78 69 79
rect 127 81 132 83
rect 127 79 128 81
rect 130 79 132 81
rect 7 72 9 74
rect 11 72 12 74
rect 7 67 12 72
rect 7 65 9 67
rect 11 65 12 67
rect 7 64 12 65
rect 7 47 11 64
rect 23 65 35 67
rect 23 63 26 65
rect 28 63 35 65
rect 23 61 35 63
rect 23 56 27 61
rect 23 54 24 56
rect 26 54 27 56
rect 23 53 27 54
rect 39 65 43 67
rect 41 63 43 65
rect 39 51 43 63
rect 47 58 51 78
rect 47 56 53 58
rect 47 54 50 56
rect 52 54 53 56
rect 47 51 53 54
rect 7 45 9 47
rect 7 43 11 45
rect 7 40 19 43
rect 7 38 9 40
rect 11 38 19 40
rect 7 37 19 38
rect 31 49 53 51
rect 31 47 50 49
rect 52 47 53 49
rect 31 45 53 47
rect 80 66 84 75
rect 127 77 132 79
rect 136 81 165 82
rect 136 79 137 81
rect 139 79 146 81
rect 148 79 165 81
rect 136 78 165 79
rect 223 81 228 83
rect 223 79 224 81
rect 226 79 228 81
rect 136 77 147 78
rect 128 72 132 77
rect 128 70 129 72
rect 131 70 132 72
rect 71 65 86 66
rect 71 63 75 65
rect 77 63 82 65
rect 84 63 86 65
rect 71 62 86 63
rect 96 65 104 67
rect 96 63 101 65
rect 103 63 104 65
rect 96 61 104 63
rect 96 58 101 61
rect 63 57 101 58
rect 63 55 64 57
rect 66 55 101 57
rect 63 54 101 55
rect 128 55 132 70
rect 127 53 132 55
rect 127 51 128 53
rect 130 51 132 53
rect 127 46 132 51
rect 127 44 128 46
rect 130 44 132 46
rect 143 58 147 77
rect 176 72 180 75
rect 176 70 177 72
rect 179 70 180 72
rect 223 77 228 79
rect 143 56 149 58
rect 143 54 146 56
rect 148 54 149 56
rect 143 49 149 54
rect 143 47 146 49
rect 148 47 149 49
rect 143 45 149 47
rect 176 66 180 70
rect 224 71 228 77
rect 224 69 225 71
rect 227 69 228 71
rect 167 65 182 66
rect 167 63 171 65
rect 173 63 178 65
rect 180 63 182 65
rect 167 62 182 63
rect 192 65 200 67
rect 192 63 197 65
rect 199 63 200 65
rect 192 62 200 63
rect 192 60 193 62
rect 195 61 200 62
rect 195 60 197 61
rect 192 58 197 60
rect 159 54 197 58
rect 224 55 228 69
rect 246 81 251 83
rect 246 79 248 81
rect 250 79 251 81
rect 246 74 251 79
rect 286 81 308 82
rect 286 79 289 81
rect 291 79 308 81
rect 286 78 308 79
rect 366 81 371 83
rect 366 79 367 81
rect 369 79 371 81
rect 246 72 248 74
rect 250 72 251 74
rect 246 70 251 72
rect 246 63 250 70
rect 232 62 250 63
rect 232 60 233 62
rect 235 60 250 62
rect 232 59 250 60
rect 223 53 228 55
rect 223 51 224 53
rect 226 51 228 53
rect 223 46 228 51
rect 127 42 132 44
rect 223 44 224 46
rect 226 44 228 46
rect 223 42 228 44
rect 119 38 132 42
rect 215 38 228 42
rect 246 47 250 59
rect 262 65 274 67
rect 262 63 265 65
rect 267 63 274 65
rect 262 61 274 63
rect 262 56 266 61
rect 262 54 263 56
rect 265 54 266 56
rect 262 53 266 54
rect 278 65 282 67
rect 280 63 282 65
rect 278 51 282 63
rect 286 58 290 78
rect 286 56 292 58
rect 286 54 289 56
rect 291 54 292 56
rect 286 51 292 54
rect 246 45 248 47
rect 246 43 250 45
rect 246 40 258 43
rect 246 38 248 40
rect 250 38 258 40
rect 246 37 258 38
rect 270 49 292 51
rect 270 47 289 49
rect 291 47 292 49
rect 270 45 292 47
rect 319 66 323 75
rect 366 77 371 79
rect 375 81 404 82
rect 375 79 376 81
rect 378 79 385 81
rect 387 79 404 81
rect 375 78 404 79
rect 462 81 467 83
rect 462 79 463 81
rect 465 79 467 81
rect 375 77 386 78
rect 367 72 371 77
rect 367 70 368 72
rect 370 70 371 72
rect 310 65 325 66
rect 310 63 314 65
rect 316 63 321 65
rect 323 63 325 65
rect 310 62 325 63
rect 335 65 343 67
rect 335 63 340 65
rect 342 63 343 65
rect 335 61 343 63
rect 335 58 340 61
rect 302 57 340 58
rect 302 55 308 57
rect 310 55 340 57
rect 302 54 340 55
rect 367 55 371 70
rect 366 53 371 55
rect 366 51 367 53
rect 369 51 371 53
rect 366 46 371 51
rect 366 44 367 46
rect 369 44 371 46
rect 382 58 386 77
rect 415 72 419 75
rect 415 70 416 72
rect 418 70 419 72
rect 462 77 467 79
rect 382 56 388 58
rect 382 54 385 56
rect 387 54 388 56
rect 382 49 388 54
rect 382 47 385 49
rect 387 47 388 49
rect 382 45 388 47
rect 415 66 419 70
rect 406 65 421 66
rect 406 63 410 65
rect 412 63 417 65
rect 419 63 421 65
rect 406 62 421 63
rect 431 65 439 67
rect 431 63 436 65
rect 438 63 439 65
rect 431 62 439 63
rect 431 60 432 62
rect 434 61 439 62
rect 434 60 436 61
rect 431 58 436 60
rect 398 54 436 58
rect 463 55 467 77
rect 462 53 467 55
rect 558 82 564 83
rect 558 80 560 82
rect 562 80 564 82
rect 558 79 564 80
rect 512 74 524 75
rect 512 72 517 74
rect 519 72 524 74
rect 512 69 524 72
rect 518 65 524 69
rect 518 63 519 65
rect 521 63 524 65
rect 518 61 524 63
rect 535 63 550 66
rect 535 61 546 63
rect 548 61 550 63
rect 535 60 550 61
rect 535 57 541 60
rect 535 55 536 57
rect 538 55 541 57
rect 535 54 541 55
rect 462 51 463 53
rect 465 51 467 53
rect 462 46 467 51
rect 560 50 564 79
rect 366 42 371 44
rect 462 44 463 46
rect 465 44 467 46
rect 462 43 467 44
rect 462 42 464 43
rect 358 38 371 42
rect 454 41 464 42
rect 466 41 467 43
rect 454 38 467 41
rect 504 47 517 50
rect 504 45 506 47
rect 508 46 517 47
rect 551 48 564 50
rect 551 46 560 48
rect 562 46 564 48
rect 508 45 509 46
rect 558 45 564 46
rect 504 37 509 45
rect 3 31 568 32
rect 3 29 20 31
rect 22 29 259 31
rect 261 29 507 31
rect 509 29 568 31
rect 3 19 568 29
rect 3 17 213 19
rect 215 17 453 19
rect 455 17 507 19
rect 509 17 568 19
rect 3 16 568 17
rect 7 6 20 10
rect 103 6 116 10
rect 7 4 12 6
rect 7 2 9 4
rect 11 2 12 4
rect 103 4 108 6
rect 7 -3 12 2
rect 7 -5 9 -3
rect 11 -5 12 -3
rect 7 -7 12 -5
rect 7 -29 11 -7
rect 38 -10 76 -6
rect 38 -13 43 -10
rect 35 -15 43 -13
rect 35 -17 36 -15
rect 38 -17 43 -15
rect 35 -19 43 -17
rect 53 -15 68 -14
rect 53 -17 55 -15
rect 57 -17 62 -15
rect 64 -17 68 -15
rect 53 -18 68 -17
rect 55 -22 59 -18
rect 86 1 92 3
rect 86 -1 87 1
rect 89 -1 92 1
rect 86 -6 92 -1
rect 86 -8 87 -6
rect 89 -8 92 -6
rect 86 -10 92 -8
rect 7 -31 12 -29
rect 55 -24 56 -22
rect 58 -24 59 -22
rect 55 -27 59 -24
rect 88 -29 92 -10
rect 103 2 105 4
rect 107 2 108 4
rect 103 -3 108 2
rect 103 -5 105 -3
rect 107 -5 108 -3
rect 103 -7 108 -5
rect 103 -22 107 -7
rect 134 -10 172 -6
rect 134 -13 139 -10
rect 131 -15 139 -13
rect 131 -17 132 -15
rect 134 -17 139 -15
rect 131 -19 139 -17
rect 149 -15 164 -14
rect 149 -17 151 -15
rect 153 -17 158 -15
rect 160 -17 164 -15
rect 149 -18 164 -17
rect 103 -24 104 -22
rect 106 -24 107 -22
rect 103 -29 107 -24
rect 88 -30 99 -29
rect 7 -33 9 -31
rect 11 -33 12 -31
rect 7 -35 12 -33
rect 70 -31 99 -30
rect 70 -33 87 -31
rect 89 -33 96 -31
rect 98 -33 99 -31
rect 70 -34 99 -33
rect 103 -31 108 -29
rect 151 -27 155 -18
rect 182 1 204 3
rect 182 -1 183 1
rect 185 -1 204 1
rect 182 -3 204 -1
rect 216 10 228 11
rect 216 8 224 10
rect 226 8 228 10
rect 216 5 228 8
rect 224 3 228 5
rect 226 1 228 3
rect 182 -6 188 -3
rect 182 -8 183 -6
rect 185 -8 188 -6
rect 182 -10 188 -8
rect 184 -30 188 -10
rect 192 -15 196 -3
rect 192 -17 194 -15
rect 192 -19 196 -17
rect 208 -6 212 -5
rect 208 -8 209 -6
rect 211 -8 212 -6
rect 208 -13 212 -8
rect 200 -15 212 -13
rect 200 -17 207 -15
rect 209 -17 212 -15
rect 200 -19 212 -17
rect 224 -11 228 1
rect 247 6 260 10
rect 343 6 356 10
rect 247 4 252 6
rect 247 2 249 4
rect 251 2 252 4
rect 343 4 348 6
rect 247 -3 252 2
rect 247 -5 249 -3
rect 251 -5 252 -3
rect 247 -7 252 -5
rect 224 -12 243 -11
rect 224 -14 240 -12
rect 242 -14 243 -12
rect 224 -15 243 -14
rect 224 -22 228 -15
rect 223 -24 228 -22
rect 223 -26 224 -24
rect 226 -26 228 -24
rect 103 -33 105 -31
rect 107 -33 108 -31
rect 103 -35 108 -33
rect 166 -31 188 -30
rect 166 -33 183 -31
rect 185 -33 188 -31
rect 166 -34 188 -33
rect 223 -31 228 -26
rect 223 -33 224 -31
rect 226 -33 228 -31
rect 223 -35 228 -33
rect 247 -29 251 -7
rect 278 -10 316 -6
rect 278 -12 283 -10
rect 278 -13 280 -12
rect 275 -14 280 -13
rect 282 -14 283 -12
rect 275 -15 283 -14
rect 275 -17 276 -15
rect 278 -17 283 -15
rect 275 -19 283 -17
rect 293 -15 308 -14
rect 293 -17 295 -15
rect 297 -17 302 -15
rect 304 -17 308 -15
rect 293 -18 308 -17
rect 295 -22 299 -18
rect 326 1 332 3
rect 326 -1 327 1
rect 329 -1 332 1
rect 326 -6 332 -1
rect 326 -8 327 -6
rect 329 -8 332 -6
rect 326 -10 332 -8
rect 247 -31 252 -29
rect 295 -24 296 -22
rect 298 -24 299 -22
rect 295 -27 299 -24
rect 328 -29 332 -10
rect 343 2 345 4
rect 347 2 348 4
rect 343 -3 348 2
rect 343 -5 345 -3
rect 347 -5 348 -3
rect 343 -7 348 -5
rect 343 -22 347 -7
rect 374 -10 412 -6
rect 374 -13 379 -10
rect 371 -15 379 -13
rect 371 -17 372 -15
rect 374 -17 379 -15
rect 371 -19 379 -17
rect 389 -15 404 -14
rect 389 -17 391 -15
rect 393 -17 398 -15
rect 400 -17 404 -15
rect 389 -18 404 -17
rect 343 -24 344 -22
rect 346 -24 347 -22
rect 343 -29 347 -24
rect 328 -30 339 -29
rect 247 -33 249 -31
rect 251 -33 252 -31
rect 247 -35 252 -33
rect 310 -31 339 -30
rect 310 -33 327 -31
rect 329 -33 336 -31
rect 338 -33 339 -31
rect 310 -34 339 -33
rect 343 -31 348 -29
rect 391 -27 395 -18
rect 422 1 444 3
rect 422 -1 423 1
rect 425 -1 444 1
rect 422 -3 444 -1
rect 456 10 468 11
rect 456 8 464 10
rect 466 8 468 10
rect 456 5 468 8
rect 464 3 468 5
rect 466 1 468 3
rect 422 -6 428 -3
rect 422 -8 423 -6
rect 425 -8 428 -6
rect 422 -10 428 -8
rect 424 -30 428 -10
rect 432 -15 436 -3
rect 432 -17 434 -15
rect 432 -19 436 -17
rect 448 -6 452 -5
rect 448 -8 449 -6
rect 451 -8 452 -6
rect 448 -13 452 -8
rect 440 -15 452 -13
rect 440 -17 447 -15
rect 449 -17 452 -15
rect 440 -19 452 -17
rect 464 -11 468 1
rect 504 3 509 11
rect 504 1 506 3
rect 508 2 509 3
rect 558 2 564 3
rect 508 1 517 2
rect 504 -2 517 1
rect 551 0 560 2
rect 562 0 564 2
rect 551 -2 564 0
rect 464 -12 484 -11
rect 464 -14 481 -12
rect 483 -14 484 -12
rect 464 -15 484 -14
rect 464 -22 468 -15
rect 463 -24 468 -22
rect 463 -26 464 -24
rect 466 -26 468 -24
rect 343 -33 345 -31
rect 347 -33 348 -31
rect 343 -35 348 -33
rect 406 -31 428 -30
rect 406 -33 423 -31
rect 425 -33 428 -31
rect 406 -34 428 -33
rect 463 -31 468 -26
rect 463 -33 464 -31
rect 466 -33 468 -31
rect 463 -35 468 -33
rect 518 -15 524 -13
rect 518 -17 519 -15
rect 521 -17 524 -15
rect 518 -21 524 -17
rect 512 -24 524 -21
rect 512 -26 517 -24
rect 519 -26 524 -24
rect 512 -27 524 -26
rect 535 -7 541 -6
rect 535 -9 536 -7
rect 538 -9 541 -7
rect 535 -12 541 -9
rect 535 -13 550 -12
rect 535 -15 546 -13
rect 548 -15 550 -13
rect 535 -18 550 -15
rect 560 -31 564 -2
rect 558 -32 564 -31
rect 558 -34 560 -32
rect 562 -34 564 -32
rect 558 -35 564 -34
rect 3 -41 568 -40
rect 3 -43 197 -41
rect 199 -43 437 -41
rect 439 -43 568 -41
rect 3 -53 568 -43
rect 3 -55 36 -53
rect 38 -55 275 -53
rect 277 -55 568 -53
rect 3 -56 568 -55
rect 7 -63 12 -61
rect 7 -65 9 -63
rect 11 -65 12 -63
rect 7 -70 12 -65
rect 47 -63 69 -62
rect 47 -65 50 -63
rect 52 -65 69 -63
rect 47 -66 69 -65
rect 127 -63 132 -61
rect 127 -65 128 -63
rect 130 -65 132 -63
rect 7 -72 9 -70
rect 11 -72 12 -70
rect 7 -74 12 -72
rect 7 -97 11 -74
rect 23 -79 35 -77
rect 23 -81 26 -79
rect 28 -81 35 -79
rect 23 -83 35 -81
rect 23 -88 27 -83
rect 23 -90 24 -88
rect 26 -90 27 -88
rect 23 -91 27 -90
rect 39 -79 43 -77
rect 41 -81 43 -79
rect 39 -93 43 -81
rect 47 -86 51 -66
rect 47 -88 53 -86
rect 47 -90 50 -88
rect 52 -90 53 -88
rect 47 -93 53 -90
rect 7 -99 9 -97
rect 7 -101 11 -99
rect 7 -104 19 -101
rect 7 -106 9 -104
rect 11 -106 19 -104
rect 7 -107 19 -106
rect 31 -95 53 -93
rect 31 -97 50 -95
rect 52 -97 53 -95
rect 31 -99 53 -97
rect 80 -78 84 -69
rect 127 -67 132 -65
rect 136 -63 165 -62
rect 136 -65 137 -63
rect 139 -65 146 -63
rect 148 -65 165 -63
rect 136 -66 165 -65
rect 223 -63 228 -61
rect 223 -65 224 -63
rect 226 -65 228 -63
rect 136 -67 147 -66
rect 128 -72 132 -67
rect 128 -74 129 -72
rect 131 -74 132 -72
rect 71 -79 86 -78
rect 71 -81 75 -79
rect 77 -81 82 -79
rect 84 -81 86 -79
rect 71 -82 86 -81
rect 96 -79 104 -77
rect 96 -81 101 -79
rect 103 -81 104 -79
rect 96 -83 104 -81
rect 96 -86 101 -83
rect 63 -87 101 -86
rect 63 -89 64 -87
rect 66 -89 101 -87
rect 63 -90 101 -89
rect 128 -89 132 -74
rect 127 -91 132 -89
rect 127 -93 128 -91
rect 130 -93 132 -91
rect 127 -98 132 -93
rect 127 -100 128 -98
rect 130 -100 132 -98
rect 143 -86 147 -67
rect 176 -72 180 -69
rect 176 -74 177 -72
rect 179 -74 180 -72
rect 223 -67 228 -65
rect 143 -88 149 -86
rect 143 -90 146 -88
rect 148 -90 149 -88
rect 143 -95 149 -90
rect 143 -97 146 -95
rect 148 -97 149 -95
rect 143 -99 149 -97
rect 176 -78 180 -74
rect 167 -79 182 -78
rect 167 -81 171 -79
rect 173 -81 178 -79
rect 180 -81 182 -79
rect 167 -82 182 -81
rect 192 -79 200 -77
rect 192 -81 197 -79
rect 199 -81 200 -79
rect 192 -82 200 -81
rect 192 -84 193 -82
rect 195 -83 200 -82
rect 195 -84 197 -83
rect 192 -86 197 -84
rect 159 -90 197 -86
rect 224 -89 228 -67
rect 246 -63 251 -61
rect 246 -65 248 -63
rect 250 -65 251 -63
rect 246 -70 251 -65
rect 286 -63 308 -62
rect 286 -65 289 -63
rect 291 -65 308 -63
rect 286 -66 308 -65
rect 366 -63 371 -61
rect 366 -65 367 -63
rect 369 -65 371 -63
rect 246 -72 248 -70
rect 250 -72 251 -70
rect 246 -74 251 -72
rect 246 -81 250 -74
rect 232 -82 250 -81
rect 232 -84 233 -82
rect 235 -84 250 -82
rect 232 -85 250 -84
rect 223 -91 228 -89
rect 223 -93 224 -91
rect 226 -93 228 -91
rect 223 -98 228 -93
rect 127 -102 132 -100
rect 223 -100 224 -98
rect 226 -100 228 -98
rect 223 -102 228 -100
rect 119 -106 132 -102
rect 215 -106 228 -102
rect 246 -97 250 -85
rect 262 -79 274 -77
rect 262 -81 265 -79
rect 267 -81 274 -79
rect 262 -83 274 -81
rect 262 -88 266 -83
rect 262 -90 263 -88
rect 265 -90 266 -88
rect 262 -91 266 -90
rect 278 -79 282 -77
rect 280 -81 282 -79
rect 278 -93 282 -81
rect 286 -86 290 -66
rect 286 -88 292 -86
rect 286 -90 289 -88
rect 291 -90 292 -88
rect 286 -93 292 -90
rect 246 -99 248 -97
rect 246 -101 250 -99
rect 246 -104 258 -101
rect 246 -106 248 -104
rect 250 -106 258 -104
rect 246 -107 258 -106
rect 270 -95 292 -93
rect 270 -97 289 -95
rect 291 -97 292 -95
rect 270 -99 292 -97
rect 319 -78 323 -69
rect 366 -67 371 -65
rect 375 -63 404 -62
rect 375 -65 376 -63
rect 378 -65 385 -63
rect 387 -65 404 -63
rect 375 -66 404 -65
rect 462 -63 467 -61
rect 462 -65 463 -63
rect 465 -65 467 -63
rect 375 -67 386 -66
rect 367 -72 371 -67
rect 367 -74 368 -72
rect 370 -74 371 -72
rect 310 -79 325 -78
rect 310 -81 314 -79
rect 316 -81 321 -79
rect 323 -81 325 -79
rect 310 -82 325 -81
rect 335 -79 343 -77
rect 335 -81 340 -79
rect 342 -81 343 -79
rect 335 -83 343 -81
rect 335 -86 340 -83
rect 302 -90 340 -86
rect 367 -89 371 -74
rect 366 -91 371 -89
rect 366 -93 367 -91
rect 369 -93 371 -91
rect 366 -98 371 -93
rect 366 -100 367 -98
rect 369 -100 371 -98
rect 382 -86 386 -67
rect 415 -72 419 -69
rect 415 -74 416 -72
rect 418 -74 419 -72
rect 462 -67 467 -65
rect 382 -88 388 -86
rect 382 -90 385 -88
rect 387 -90 388 -88
rect 382 -95 388 -90
rect 382 -97 385 -95
rect 387 -97 388 -95
rect 382 -99 388 -97
rect 415 -78 419 -74
rect 406 -79 421 -78
rect 406 -81 410 -79
rect 412 -81 417 -79
rect 419 -81 421 -79
rect 406 -82 421 -81
rect 431 -79 439 -77
rect 431 -81 436 -79
rect 438 -81 439 -79
rect 431 -82 439 -81
rect 431 -84 432 -82
rect 434 -83 439 -82
rect 434 -84 436 -83
rect 431 -86 436 -84
rect 398 -90 436 -86
rect 463 -89 467 -67
rect 462 -91 467 -89
rect 558 -62 564 -61
rect 558 -64 560 -62
rect 562 -64 564 -62
rect 558 -65 564 -64
rect 512 -75 524 -69
rect 518 -79 524 -75
rect 518 -81 519 -79
rect 521 -81 524 -79
rect 518 -83 524 -81
rect 535 -81 550 -78
rect 535 -83 546 -81
rect 548 -83 550 -81
rect 535 -84 550 -83
rect 535 -86 536 -84
rect 538 -86 541 -84
rect 535 -90 541 -86
rect 462 -93 463 -91
rect 465 -93 467 -91
rect 462 -98 467 -93
rect 560 -94 564 -65
rect 366 -102 371 -100
rect 462 -100 463 -98
rect 465 -100 467 -98
rect 462 -102 467 -100
rect 358 -106 371 -102
rect 454 -106 467 -102
rect 504 -97 517 -94
rect 504 -99 506 -97
rect 508 -98 517 -97
rect 551 -96 564 -94
rect 551 -98 560 -96
rect 562 -98 564 -96
rect 508 -99 509 -98
rect 558 -99 564 -98
rect 504 -107 509 -99
rect 3 -113 568 -112
rect 3 -115 20 -113
rect 22 -115 259 -113
rect 261 -115 507 -113
rect 509 -115 568 -113
rect 3 -120 568 -115
<< alu2 >>
rect 87 217 91 218
rect 87 215 88 217
rect 90 215 91 217
rect 87 214 91 215
rect 88 209 92 210
rect 88 207 89 209
rect 91 207 92 209
rect 88 206 92 207
rect 24 205 28 206
rect 24 203 25 205
rect 27 203 28 205
rect 24 202 28 203
rect 245 201 249 202
rect 245 199 246 201
rect 248 199 249 201
rect 245 198 249 199
rect 307 201 358 202
rect 307 199 308 201
rect 310 199 354 201
rect 356 199 358 201
rect 307 198 358 199
rect 196 195 200 196
rect 116 193 120 194
rect 196 193 197 195
rect 199 193 200 195
rect 63 192 67 193
rect 63 190 64 192
rect 66 190 67 192
rect 116 191 117 193
rect 119 191 120 193
rect 116 190 120 191
rect 142 192 146 193
rect 196 192 200 193
rect 422 193 426 194
rect 142 190 143 192
rect 145 190 146 192
rect 422 191 423 193
rect 425 191 426 193
rect 422 190 426 191
rect 474 193 478 194
rect 474 191 475 193
rect 477 191 478 193
rect 474 190 478 191
rect 516 193 520 194
rect 516 191 517 193
rect 519 191 520 193
rect 516 190 520 191
rect 560 193 564 194
rect 560 191 561 193
rect 563 191 564 193
rect 560 190 564 191
rect 63 189 67 190
rect 142 189 146 190
rect 96 184 100 185
rect 96 182 97 184
rect 99 182 100 184
rect 96 181 100 182
rect 128 184 132 185
rect 128 182 129 184
rect 131 182 132 184
rect 128 181 132 182
rect 212 184 216 185
rect 212 182 213 184
rect 215 182 216 184
rect 212 181 216 182
rect 322 184 327 185
rect 322 182 323 184
rect 325 182 327 184
rect 322 181 327 182
rect 7 153 11 154
rect 7 151 8 153
rect 10 151 11 153
rect 7 150 11 151
rect 208 138 234 139
rect 448 138 474 139
rect 150 137 154 138
rect 150 135 151 137
rect 153 135 154 137
rect 150 134 154 135
rect 208 136 209 138
rect 211 136 234 138
rect 208 134 234 136
rect 375 137 379 138
rect 375 135 376 137
rect 378 135 379 137
rect 375 134 379 135
rect 448 136 449 138
rect 451 136 474 138
rect 448 134 474 136
rect 55 122 107 123
rect 55 120 56 122
rect 58 120 104 122
rect 106 120 107 122
rect 55 119 107 120
rect 230 115 234 134
rect 239 132 283 133
rect 239 130 240 132
rect 242 130 280 132
rect 282 130 283 132
rect 239 129 283 130
rect 247 124 251 125
rect 247 122 248 124
rect 250 122 251 124
rect 247 121 251 122
rect 295 122 347 123
rect 295 120 296 122
rect 298 120 344 122
rect 346 120 347 122
rect 295 119 347 120
rect 470 115 474 134
rect 95 113 234 115
rect 95 111 96 113
rect 98 111 234 113
rect 95 110 234 111
rect 335 113 474 115
rect 335 111 336 113
rect 338 111 474 113
rect 335 110 474 111
rect 480 132 485 133
rect 480 130 481 132
rect 483 130 485 132
rect 0 81 140 82
rect 0 79 137 81
rect 139 79 140 81
rect 0 77 140 79
rect 240 81 379 82
rect 240 79 376 81
rect 378 79 379 81
rect 240 77 379 79
rect 0 58 4 77
rect 128 72 180 73
rect 128 70 129 72
rect 131 70 177 72
rect 179 70 180 72
rect 128 69 180 70
rect 224 71 228 72
rect 224 69 225 71
rect 227 69 228 71
rect 224 68 228 69
rect 8 67 12 68
rect 8 65 9 67
rect 11 65 12 67
rect 8 64 12 65
rect 192 62 236 63
rect 192 60 193 62
rect 195 60 233 62
rect 235 60 236 62
rect 192 59 236 60
rect 240 58 244 77
rect 367 72 419 73
rect 367 70 368 72
rect 370 70 416 72
rect 418 70 419 72
rect 367 69 419 70
rect 480 63 485 130
rect 513 122 517 123
rect 513 120 514 122
rect 516 120 517 122
rect 513 119 517 120
rect 516 74 520 75
rect 516 72 517 74
rect 519 72 520 74
rect 516 71 520 72
rect 431 62 485 63
rect 431 60 432 62
rect 434 60 485 62
rect 431 59 485 60
rect 0 56 27 58
rect 0 54 24 56
rect 26 54 27 56
rect 63 57 67 58
rect 63 55 64 57
rect 66 55 67 57
rect 63 54 67 55
rect 240 56 266 58
rect 240 54 263 56
rect 265 54 266 56
rect 307 57 311 58
rect 307 55 308 57
rect 310 55 311 57
rect 307 54 311 55
rect 535 57 539 58
rect 535 55 536 57
rect 538 55 539 57
rect 535 54 539 55
rect 0 53 27 54
rect 240 53 266 54
rect 463 43 467 44
rect 463 41 464 43
rect 466 41 467 43
rect 463 40 467 41
rect 208 -6 234 -5
rect 208 -8 209 -6
rect 211 -8 234 -6
rect 208 -10 234 -8
rect 448 -6 474 -5
rect 448 -8 449 -6
rect 451 -8 474 -6
rect 448 -10 474 -8
rect 535 -7 539 -6
rect 535 -9 536 -7
rect 538 -9 539 -7
rect 535 -10 539 -9
rect 55 -22 107 -21
rect 55 -24 56 -22
rect 58 -24 104 -22
rect 106 -24 107 -22
rect 55 -25 107 -24
rect 230 -29 234 -10
rect 239 -12 283 -11
rect 239 -14 240 -12
rect 242 -14 280 -12
rect 282 -14 283 -12
rect 239 -15 283 -14
rect 295 -22 347 -21
rect 295 -24 296 -22
rect 298 -24 344 -22
rect 346 -24 347 -22
rect 295 -25 347 -24
rect 470 -29 474 -10
rect 95 -31 234 -29
rect 95 -33 96 -31
rect 98 -33 234 -31
rect 95 -34 234 -33
rect 335 -31 474 -29
rect 335 -33 336 -31
rect 338 -33 474 -31
rect 335 -34 474 -33
rect 480 -12 485 -11
rect 480 -14 481 -12
rect 483 -14 485 -12
rect 1 -63 140 -62
rect 1 -65 137 -63
rect 139 -65 140 -63
rect 1 -67 140 -65
rect 240 -63 379 -62
rect 240 -65 376 -63
rect 378 -65 379 -63
rect 240 -67 379 -65
rect 1 -86 5 -67
rect 128 -72 180 -71
rect 128 -74 129 -72
rect 131 -74 177 -72
rect 179 -74 180 -72
rect 128 -75 180 -74
rect 192 -82 236 -81
rect 192 -84 193 -82
rect 195 -84 233 -82
rect 235 -84 236 -82
rect 192 -85 236 -84
rect 240 -86 244 -67
rect 367 -72 419 -71
rect 367 -74 368 -72
rect 370 -74 416 -72
rect 418 -74 419 -72
rect 367 -75 419 -74
rect 480 -81 485 -14
rect 516 -24 520 -23
rect 516 -26 517 -24
rect 519 -26 520 -24
rect 516 -27 520 -26
rect 431 -82 485 -81
rect 431 -84 432 -82
rect 434 -84 485 -82
rect 431 -85 485 -84
rect 535 -84 539 -83
rect 535 -86 536 -84
rect 538 -86 539 -84
rect 1 -88 27 -86
rect 1 -90 24 -88
rect 26 -90 27 -88
rect 63 -87 67 -86
rect 63 -89 64 -87
rect 66 -89 67 -87
rect 63 -90 67 -89
rect 240 -88 266 -86
rect 535 -87 539 -86
rect 240 -90 263 -88
rect 265 -90 266 -88
rect 1 -91 27 -90
rect 240 -91 266 -90
<< alu3 >>
rect 7 217 91 218
rect 7 215 8 217
rect 10 215 88 217
rect 90 215 91 217
rect 7 214 91 215
rect 88 209 92 210
rect 88 207 89 209
rect 91 207 92 209
rect 88 206 92 207
rect 24 205 28 206
rect 24 203 25 205
rect 27 203 28 205
rect 24 202 28 203
rect 245 201 249 202
rect 245 199 246 201
rect 248 199 249 201
rect 245 198 249 199
rect 196 195 200 196
rect 116 193 120 194
rect 196 193 197 195
rect 199 193 200 195
rect 63 192 67 193
rect 63 190 64 192
rect 66 190 67 192
rect 116 191 117 193
rect 119 191 120 193
rect 116 190 120 191
rect 142 192 146 193
rect 196 192 200 193
rect 422 193 426 194
rect 142 190 143 192
rect 145 190 146 192
rect 422 191 423 193
rect 425 191 426 193
rect 422 190 426 191
rect 474 193 478 194
rect 474 191 475 193
rect 477 191 478 193
rect 474 190 478 191
rect 516 193 520 194
rect 516 191 517 193
rect 519 191 520 193
rect 516 190 520 191
rect 560 193 564 194
rect 560 191 561 193
rect 563 191 564 193
rect 560 190 564 191
rect 63 189 67 190
rect 142 189 146 190
rect 96 184 100 185
rect 96 182 97 184
rect 99 182 100 184
rect 96 181 100 182
rect 128 184 327 185
rect 128 182 129 184
rect 131 182 213 184
rect 215 182 323 184
rect 325 182 327 184
rect 128 181 327 182
rect 24 165 154 166
rect 24 163 25 165
rect 27 163 151 165
rect 153 163 154 165
rect 24 162 154 163
rect 7 153 11 154
rect 7 151 8 153
rect 10 151 11 153
rect 7 150 11 151
rect 150 137 154 138
rect 150 135 151 137
rect 153 135 154 137
rect 150 134 154 135
rect 196 137 379 138
rect 196 135 197 137
rect 199 135 376 137
rect 378 135 379 137
rect 196 134 379 135
rect 116 127 251 128
rect 116 125 117 127
rect 119 125 251 127
rect 116 124 251 125
rect 247 122 248 124
rect 250 122 251 124
rect 247 121 251 122
rect 474 122 517 123
rect 474 120 475 122
rect 477 120 514 122
rect 516 120 517 122
rect 474 119 517 120
rect 516 74 520 75
rect 516 72 517 74
rect 519 72 520 74
rect 88 71 228 72
rect 516 71 520 72
rect 88 69 89 71
rect 91 69 225 71
rect 227 69 228 71
rect 88 68 228 69
rect 8 67 12 68
rect 8 65 9 67
rect 11 65 12 67
rect 8 64 12 65
rect 63 57 67 58
rect 63 55 64 57
rect 66 55 67 57
rect 63 54 67 55
rect 142 57 311 58
rect 142 55 143 57
rect 145 55 308 57
rect 310 55 311 57
rect 142 54 311 55
rect 422 57 539 58
rect 422 55 423 57
rect 425 55 536 57
rect 538 55 539 57
rect 422 54 539 55
rect 96 43 467 44
rect 96 41 97 43
rect 99 41 464 43
rect 466 41 467 43
rect 96 40 467 41
rect 24 21 154 22
rect 24 19 25 21
rect 27 19 151 21
rect 153 19 154 21
rect 24 18 154 19
rect 474 -7 539 -6
rect 474 -9 475 -7
rect 477 -9 536 -7
rect 538 -9 539 -7
rect 474 -10 539 -9
rect 516 -24 564 -23
rect 516 -26 517 -24
rect 519 -26 561 -24
rect 563 -26 564 -24
rect 516 -27 564 -26
rect 516 -84 539 -83
rect 516 -86 517 -84
rect 519 -86 536 -84
rect 538 -86 539 -84
rect 63 -87 67 -86
rect 516 -87 539 -86
rect 63 -89 64 -87
rect 66 -89 67 -87
rect 63 -90 67 -89
<< alu4 >>
rect 7 217 11 218
rect 7 215 8 217
rect 10 215 11 217
rect 7 153 11 215
rect 88 209 92 210
rect 88 207 89 209
rect 91 207 92 209
rect 24 205 28 206
rect 24 203 25 205
rect 27 203 28 205
rect 24 165 28 203
rect 24 163 25 165
rect 27 163 28 165
rect 24 162 28 163
rect 63 192 67 193
rect 63 190 64 192
rect 66 190 67 192
rect 7 151 8 153
rect 10 151 11 153
rect 7 150 11 151
rect 8 67 12 68
rect 8 65 9 67
rect 11 65 12 67
rect 8 64 12 65
rect 63 57 67 190
rect 88 71 92 207
rect 245 201 249 202
rect 245 199 246 201
rect 248 199 249 201
rect 196 195 200 197
rect 116 193 120 194
rect 196 193 197 195
rect 199 193 200 195
rect 116 191 117 193
rect 119 191 120 193
rect 88 69 89 71
rect 91 69 92 71
rect 88 68 92 69
rect 96 184 100 185
rect 96 182 97 184
rect 99 182 100 184
rect 63 55 64 57
rect 66 55 67 57
rect 63 54 67 55
rect 96 43 100 182
rect 116 127 120 191
rect 116 125 117 127
rect 119 125 120 127
rect 116 124 120 125
rect 142 192 146 193
rect 142 190 143 192
rect 145 190 146 192
rect 142 57 146 190
rect 150 165 154 166
rect 150 163 151 165
rect 153 163 154 165
rect 150 137 154 163
rect 150 135 151 137
rect 153 135 154 137
rect 150 134 154 135
rect 196 137 200 193
rect 196 135 197 137
rect 199 135 200 137
rect 196 134 200 135
rect 245 67 249 199
rect 245 65 246 67
rect 248 65 249 67
rect 245 64 249 65
rect 422 193 426 194
rect 422 191 423 193
rect 425 191 426 193
rect 142 55 143 57
rect 145 55 146 57
rect 142 54 146 55
rect 422 57 426 191
rect 422 55 423 57
rect 425 55 426 57
rect 422 54 426 55
rect 474 193 478 194
rect 474 191 475 193
rect 477 191 478 193
rect 474 122 478 191
rect 474 120 475 122
rect 477 120 478 122
rect 96 41 97 43
rect 99 41 100 43
rect 96 40 100 41
rect 24 21 28 24
rect 24 19 25 21
rect 27 19 28 21
rect 24 18 28 19
rect 63 -87 67 24
rect 150 21 154 22
rect 150 19 151 21
rect 153 19 154 21
rect 150 -6 154 19
rect 474 -7 478 120
rect 474 -9 475 -7
rect 477 -9 478 -7
rect 474 -10 478 -9
rect 516 193 520 194
rect 516 191 517 193
rect 519 191 520 193
rect 516 74 520 191
rect 516 72 517 74
rect 519 72 520 74
rect 516 -84 520 72
rect 560 193 564 194
rect 560 191 561 193
rect 563 191 564 193
rect 560 -24 564 191
rect 560 -26 561 -24
rect 563 -26 564 -24
rect 560 -27 564 -26
rect 516 -86 517 -84
rect 519 -86 520 -84
rect 516 -87 520 -86
rect 63 -89 64 -87
rect 66 -89 67 -87
rect 63 -90 67 -89
<< alu5 >>
rect 8 67 249 68
rect 8 65 9 67
rect 11 65 246 67
rect 248 65 249 67
rect 8 64 249 65
<< ptie >>
rect 117 235 131 237
rect 117 233 119 235
rect 121 233 127 235
rect 129 233 131 235
rect 117 231 131 233
rect 284 235 290 237
rect 284 233 286 235
rect 288 233 290 235
rect 284 231 290 233
rect 193 103 203 105
rect 193 101 197 103
rect 199 101 203 103
rect 193 99 203 101
rect 433 103 443 105
rect 433 101 437 103
rect 439 101 443 103
rect 433 99 443 101
rect 32 91 42 93
rect 32 89 36 91
rect 38 89 42 91
rect 32 87 42 89
rect 271 91 281 93
rect 271 89 275 91
rect 277 89 281 91
rect 271 87 281 89
rect 193 -41 203 -39
rect 193 -43 197 -41
rect 199 -43 203 -41
rect 193 -45 203 -43
rect 433 -41 443 -39
rect 433 -43 437 -41
rect 439 -43 443 -41
rect 433 -45 443 -43
rect 32 -53 42 -51
rect 32 -55 36 -53
rect 38 -55 42 -53
rect 32 -57 42 -55
rect 271 -53 281 -51
rect 271 -55 275 -53
rect 277 -55 281 -53
rect 271 -57 281 -55
<< ntie >>
rect 125 175 131 177
rect 125 173 127 175
rect 129 173 131 175
rect 213 175 219 177
rect 125 171 131 173
rect 213 173 215 175
rect 217 173 219 175
rect 323 175 329 177
rect 213 171 219 173
rect 323 173 325 175
rect 327 173 329 175
rect 323 171 329 173
rect 505 163 511 165
rect 505 161 507 163
rect 509 161 511 163
rect 505 159 511 161
rect 505 31 511 33
rect 505 29 507 31
rect 509 29 511 31
rect 505 27 511 29
rect 505 19 511 21
rect 505 17 507 19
rect 509 17 511 19
rect 505 15 511 17
rect 505 -113 511 -111
rect 505 -115 507 -113
rect 509 -115 511 -113
rect 505 -117 511 -115
<< nmos >>
rect 19 214 21 228
rect 52 214 54 228
rect 93 221 95 227
rect 103 221 105 227
rect 113 219 115 225
rect 123 219 125 225
rect 153 214 155 228
rect 189 214 191 228
rect 219 222 221 228
rect 229 222 231 228
rect 236 222 238 228
rect 246 222 248 228
rect 253 222 255 228
rect 263 222 265 228
rect 292 214 294 225
rect 302 214 304 231
rect 329 222 331 228
rect 339 222 341 228
rect 346 222 348 228
rect 356 222 358 228
rect 363 222 365 228
rect 373 222 375 228
rect 397 215 399 229
rect 407 215 409 229
rect 417 215 419 229
rect 449 215 451 229
rect 459 215 461 229
rect 469 215 471 229
rect 491 215 493 229
rect 501 215 503 229
rect 511 215 513 229
rect 535 215 537 229
rect 545 215 547 229
rect 555 215 557 229
rect 14 102 16 115
rect 24 105 26 115
rect 34 108 36 122
rect 44 108 46 122
rect 64 102 66 122
rect 71 102 73 122
rect 82 102 84 116
rect 110 102 112 115
rect 120 105 122 115
rect 130 108 132 122
rect 140 108 142 122
rect 160 102 162 122
rect 167 102 169 122
rect 178 102 180 116
rect 199 111 201 119
rect 209 109 211 117
rect 219 108 221 122
rect 254 102 256 115
rect 264 105 266 115
rect 274 108 276 122
rect 284 108 286 122
rect 304 102 306 122
rect 311 102 313 122
rect 322 102 324 116
rect 350 102 352 115
rect 360 105 362 115
rect 370 108 372 122
rect 380 108 382 122
rect 400 102 402 122
rect 407 102 409 122
rect 418 102 420 116
rect 439 111 441 119
rect 449 109 451 117
rect 459 108 461 122
rect 511 108 513 114
rect 521 108 523 114
rect 528 108 530 114
rect 538 108 540 114
rect 545 108 547 114
rect 555 108 557 114
rect 14 70 16 84
rect 24 75 26 83
rect 34 73 36 81
rect 55 76 57 90
rect 66 70 68 90
rect 73 70 75 90
rect 93 70 95 84
rect 103 70 105 84
rect 113 77 115 87
rect 123 77 125 90
rect 151 76 153 90
rect 162 70 164 90
rect 169 70 171 90
rect 189 70 191 84
rect 199 70 201 84
rect 209 77 211 87
rect 219 77 221 90
rect 253 70 255 84
rect 263 75 265 83
rect 273 73 275 81
rect 294 76 296 90
rect 305 70 307 90
rect 312 70 314 90
rect 332 70 334 84
rect 342 70 344 84
rect 352 77 354 87
rect 362 77 364 90
rect 390 76 392 90
rect 401 70 403 90
rect 408 70 410 90
rect 428 70 430 84
rect 438 70 440 84
rect 448 77 450 87
rect 458 77 460 90
rect 511 78 513 84
rect 521 78 523 84
rect 528 78 530 84
rect 538 78 540 84
rect 545 78 547 84
rect 555 78 557 84
rect 14 -42 16 -29
rect 24 -39 26 -29
rect 34 -36 36 -22
rect 44 -36 46 -22
rect 64 -42 66 -22
rect 71 -42 73 -22
rect 82 -42 84 -28
rect 110 -42 112 -29
rect 120 -39 122 -29
rect 130 -36 132 -22
rect 140 -36 142 -22
rect 160 -42 162 -22
rect 167 -42 169 -22
rect 178 -42 180 -28
rect 199 -33 201 -25
rect 209 -35 211 -27
rect 219 -36 221 -22
rect 254 -42 256 -29
rect 264 -39 266 -29
rect 274 -36 276 -22
rect 284 -36 286 -22
rect 304 -42 306 -22
rect 311 -42 313 -22
rect 322 -42 324 -28
rect 350 -42 352 -29
rect 360 -39 362 -29
rect 370 -36 372 -22
rect 380 -36 382 -22
rect 400 -42 402 -22
rect 407 -42 409 -22
rect 418 -42 420 -28
rect 439 -33 441 -25
rect 449 -35 451 -27
rect 459 -36 461 -22
rect 511 -36 513 -30
rect 521 -36 523 -30
rect 528 -36 530 -30
rect 538 -36 540 -30
rect 545 -36 547 -30
rect 555 -36 557 -30
rect 14 -74 16 -60
rect 24 -69 26 -61
rect 34 -71 36 -63
rect 55 -68 57 -54
rect 66 -74 68 -54
rect 73 -74 75 -54
rect 93 -74 95 -60
rect 103 -74 105 -60
rect 113 -67 115 -57
rect 123 -67 125 -54
rect 151 -68 153 -54
rect 162 -74 164 -54
rect 169 -74 171 -54
rect 189 -74 191 -60
rect 199 -74 201 -60
rect 209 -67 211 -57
rect 219 -67 221 -54
rect 253 -74 255 -60
rect 263 -69 265 -61
rect 273 -71 275 -63
rect 294 -68 296 -54
rect 305 -74 307 -54
rect 312 -74 314 -54
rect 332 -74 334 -60
rect 342 -74 344 -60
rect 352 -67 354 -57
rect 362 -67 364 -54
rect 390 -68 392 -54
rect 401 -74 403 -54
rect 408 -74 410 -54
rect 428 -74 430 -60
rect 438 -74 440 -60
rect 448 -67 450 -57
rect 458 -67 460 -54
rect 511 -66 513 -60
rect 521 -66 523 -60
rect 528 -66 530 -60
rect 538 -66 540 -60
rect 545 -66 547 -60
rect 555 -66 557 -60
<< pmos >>
rect 19 174 21 202
rect 52 174 54 202
rect 93 174 95 196
rect 100 174 102 196
rect 107 174 109 196
rect 114 174 116 196
rect 153 174 155 202
rect 189 174 191 202
rect 219 196 221 202
rect 229 182 231 194
rect 236 182 238 194
rect 246 182 248 194
rect 253 182 255 194
rect 263 182 265 194
rect 292 174 294 202
rect 302 174 304 202
rect 329 196 331 202
rect 339 182 341 194
rect 346 182 348 194
rect 356 182 358 194
rect 363 182 365 194
rect 373 182 375 194
rect 397 174 399 202
rect 407 174 409 202
rect 417 174 419 202
rect 449 174 451 202
rect 459 174 461 202
rect 469 174 471 202
rect 491 174 493 202
rect 501 174 503 202
rect 511 174 513 202
rect 535 174 537 202
rect 545 174 547 202
rect 555 174 557 202
rect 14 137 16 162
rect 27 137 29 150
rect 37 134 39 159
rect 44 134 46 159
rect 62 134 64 162
rect 72 134 74 162
rect 82 134 84 162
rect 110 137 112 162
rect 123 137 125 150
rect 133 134 135 159
rect 140 134 142 159
rect 158 134 160 162
rect 168 134 170 162
rect 178 134 180 162
rect 199 134 201 162
rect 206 134 208 162
rect 219 134 221 162
rect 254 137 256 162
rect 267 137 269 150
rect 277 134 279 159
rect 284 134 286 159
rect 302 134 304 162
rect 312 134 314 162
rect 322 134 324 162
rect 350 137 352 162
rect 363 137 365 150
rect 373 134 375 159
rect 380 134 382 159
rect 398 134 400 162
rect 408 134 410 162
rect 418 134 420 162
rect 439 134 441 162
rect 446 134 448 162
rect 459 134 461 162
rect 521 142 523 154
rect 528 142 530 154
rect 538 142 540 154
rect 545 142 547 154
rect 555 142 557 154
rect 511 134 513 140
rect 14 30 16 58
rect 27 30 29 58
rect 34 30 36 58
rect 55 30 57 58
rect 65 30 67 58
rect 75 30 77 58
rect 93 33 95 58
rect 100 33 102 58
rect 110 42 112 55
rect 123 30 125 55
rect 151 30 153 58
rect 161 30 163 58
rect 171 30 173 58
rect 189 33 191 58
rect 196 33 198 58
rect 206 42 208 55
rect 219 30 221 55
rect 253 30 255 58
rect 266 30 268 58
rect 273 30 275 58
rect 294 30 296 58
rect 304 30 306 58
rect 314 30 316 58
rect 332 33 334 58
rect 339 33 341 58
rect 349 42 351 55
rect 362 30 364 55
rect 390 30 392 58
rect 400 30 402 58
rect 410 30 412 58
rect 428 33 430 58
rect 435 33 437 58
rect 445 42 447 55
rect 458 30 460 55
rect 511 52 513 58
rect 521 38 523 50
rect 528 38 530 50
rect 538 38 540 50
rect 545 38 547 50
rect 555 38 557 50
rect 14 -7 16 18
rect 27 -7 29 6
rect 37 -10 39 15
rect 44 -10 46 15
rect 62 -10 64 18
rect 72 -10 74 18
rect 82 -10 84 18
rect 110 -7 112 18
rect 123 -7 125 6
rect 133 -10 135 15
rect 140 -10 142 15
rect 158 -10 160 18
rect 168 -10 170 18
rect 178 -10 180 18
rect 199 -10 201 18
rect 206 -10 208 18
rect 219 -10 221 18
rect 254 -7 256 18
rect 267 -7 269 6
rect 277 -10 279 15
rect 284 -10 286 15
rect 302 -10 304 18
rect 312 -10 314 18
rect 322 -10 324 18
rect 350 -7 352 18
rect 363 -7 365 6
rect 373 -10 375 15
rect 380 -10 382 15
rect 398 -10 400 18
rect 408 -10 410 18
rect 418 -10 420 18
rect 439 -10 441 18
rect 446 -10 448 18
rect 459 -10 461 18
rect 521 -2 523 10
rect 528 -2 530 10
rect 538 -2 540 10
rect 545 -2 547 10
rect 555 -2 557 10
rect 511 -10 513 -4
rect 14 -114 16 -86
rect 27 -114 29 -86
rect 34 -114 36 -86
rect 55 -114 57 -86
rect 65 -114 67 -86
rect 75 -114 77 -86
rect 93 -111 95 -86
rect 100 -111 102 -86
rect 110 -102 112 -89
rect 123 -114 125 -89
rect 151 -114 153 -86
rect 161 -114 163 -86
rect 171 -114 173 -86
rect 189 -111 191 -86
rect 196 -111 198 -86
rect 206 -102 208 -89
rect 219 -114 221 -89
rect 253 -114 255 -86
rect 266 -114 268 -86
rect 273 -114 275 -86
rect 294 -114 296 -86
rect 304 -114 306 -86
rect 314 -114 316 -86
rect 332 -111 334 -86
rect 339 -111 341 -86
rect 349 -102 351 -89
rect 362 -114 364 -89
rect 390 -114 392 -86
rect 400 -114 402 -86
rect 410 -114 412 -86
rect 428 -111 430 -86
rect 435 -111 437 -86
rect 445 -102 447 -89
rect 458 -114 460 -89
rect 511 -92 513 -86
rect 521 -106 523 -94
rect 528 -106 530 -94
rect 538 -106 540 -94
rect 545 -106 547 -94
rect 555 -106 557 -94
<< polyct0 >>
rect 111 207 113 209
rect 244 215 246 217
rect 262 215 264 217
rect 237 199 239 201
rect 354 215 356 217
rect 372 215 374 217
rect 347 199 349 201
rect 408 208 410 210
rect 460 208 462 210
rect 502 208 504 210
rect 546 208 548 210
rect 22 130 24 132
rect 16 120 18 122
rect 72 127 74 129
rect 82 127 84 129
rect 118 130 120 132
rect 112 120 114 122
rect 168 127 170 129
rect 178 127 180 129
rect 217 127 219 129
rect 262 130 264 132
rect 256 120 258 122
rect 312 127 314 129
rect 322 127 324 129
rect 358 130 360 132
rect 352 120 354 122
rect 408 127 410 129
rect 418 127 420 129
rect 457 127 459 129
rect 529 135 531 137
rect 536 119 538 121
rect 554 119 556 121
rect 16 63 18 65
rect 55 63 57 65
rect 65 63 67 65
rect 121 70 123 72
rect 115 60 117 62
rect 151 63 153 65
rect 161 63 163 65
rect 217 70 219 72
rect 211 60 213 62
rect 255 63 257 65
rect 294 63 296 65
rect 304 63 306 65
rect 360 70 362 72
rect 354 60 356 62
rect 390 63 392 65
rect 400 63 402 65
rect 456 70 458 72
rect 450 60 452 62
rect 536 71 538 73
rect 554 71 556 73
rect 529 55 531 57
rect 22 -14 24 -12
rect 16 -24 18 -22
rect 72 -17 74 -15
rect 82 -17 84 -15
rect 118 -14 120 -12
rect 112 -24 114 -22
rect 168 -17 170 -15
rect 178 -17 180 -15
rect 217 -17 219 -15
rect 262 -14 264 -12
rect 256 -24 258 -22
rect 312 -17 314 -15
rect 322 -17 324 -15
rect 358 -14 360 -12
rect 352 -24 354 -22
rect 408 -17 410 -15
rect 418 -17 420 -15
rect 457 -17 459 -15
rect 529 -9 531 -7
rect 536 -25 538 -23
rect 554 -25 556 -23
rect 16 -81 18 -79
rect 55 -81 57 -79
rect 65 -81 67 -79
rect 121 -74 123 -72
rect 115 -84 117 -82
rect 151 -81 153 -79
rect 161 -81 163 -79
rect 217 -74 219 -72
rect 211 -84 213 -82
rect 255 -81 257 -79
rect 294 -81 296 -79
rect 304 -81 306 -79
rect 360 -74 362 -72
rect 354 -84 356 -82
rect 390 -81 392 -79
rect 400 -81 402 -79
rect 456 -74 458 -72
rect 450 -84 452 -82
rect 536 -73 538 -71
rect 554 -73 556 -71
rect 529 -89 531 -87
<< polyct1 >>
rect 16 207 18 209
rect 49 207 51 209
rect 101 214 103 216
rect 89 201 91 203
rect 121 201 123 203
rect 156 207 158 209
rect 186 207 188 209
rect 227 207 229 209
rect 254 205 256 207
rect 293 207 295 209
rect 337 207 339 209
rect 214 189 216 191
rect 364 205 366 207
rect 398 207 400 209
rect 450 207 452 209
rect 492 207 494 209
rect 536 207 538 209
rect 324 189 326 191
rect 36 127 38 129
rect 55 127 57 129
rect 62 127 64 129
rect 132 127 134 129
rect 151 127 153 129
rect 158 127 160 129
rect 194 127 196 129
rect 207 127 209 129
rect 276 127 278 129
rect 295 127 297 129
rect 302 127 304 129
rect 506 145 508 147
rect 372 127 374 129
rect 391 127 393 129
rect 398 127 400 129
rect 434 127 436 129
rect 447 127 449 129
rect 519 127 521 129
rect 546 129 548 131
rect 26 63 28 65
rect 39 63 41 65
rect 75 63 77 65
rect 82 63 84 65
rect 101 63 103 65
rect 171 63 173 65
rect 178 63 180 65
rect 197 63 199 65
rect 265 63 267 65
rect 278 63 280 65
rect 314 63 316 65
rect 321 63 323 65
rect 340 63 342 65
rect 410 63 412 65
rect 417 63 419 65
rect 436 63 438 65
rect 519 63 521 65
rect 546 61 548 63
rect 506 45 508 47
rect 36 -17 38 -15
rect 55 -17 57 -15
rect 62 -17 64 -15
rect 132 -17 134 -15
rect 151 -17 153 -15
rect 158 -17 160 -15
rect 194 -17 196 -15
rect 207 -17 209 -15
rect 276 -17 278 -15
rect 295 -17 297 -15
rect 302 -17 304 -15
rect 506 1 508 3
rect 372 -17 374 -15
rect 391 -17 393 -15
rect 398 -17 400 -15
rect 434 -17 436 -15
rect 447 -17 449 -15
rect 519 -17 521 -15
rect 546 -15 548 -13
rect 26 -81 28 -79
rect 39 -81 41 -79
rect 75 -81 77 -79
rect 82 -81 84 -79
rect 101 -81 103 -79
rect 171 -81 173 -79
rect 178 -81 180 -79
rect 197 -81 199 -79
rect 265 -81 267 -79
rect 278 -81 280 -79
rect 314 -81 316 -79
rect 321 -81 323 -79
rect 340 -81 342 -79
rect 410 -81 412 -79
rect 417 -81 419 -79
rect 436 -81 438 -79
rect 519 -81 521 -79
rect 546 -83 548 -81
rect 506 -99 508 -97
<< ndifct0 >>
rect 14 224 16 226
rect 14 217 16 219
rect 47 224 49 226
rect 47 217 49 219
rect 128 221 130 223
rect 158 224 160 226
rect 158 217 160 219
rect 184 224 186 226
rect 184 217 186 219
rect 214 224 216 226
rect 224 224 226 226
rect 241 224 243 226
rect 258 224 260 226
rect 287 220 289 222
rect 307 227 309 229
rect 324 224 326 226
rect 334 224 336 226
rect 351 224 353 226
rect 368 224 370 226
rect 392 224 394 226
rect 392 217 394 219
rect 402 225 404 227
rect 422 225 424 227
rect 422 217 424 219
rect 444 224 446 226
rect 444 217 446 219
rect 454 225 456 227
rect 474 225 476 227
rect 474 217 476 219
rect 486 224 488 226
rect 486 217 488 219
rect 496 225 498 227
rect 516 225 518 227
rect 516 217 518 219
rect 530 224 532 226
rect 530 217 532 219
rect 540 225 542 227
rect 560 225 562 227
rect 560 217 562 219
rect 19 107 21 109
rect 29 110 31 112
rect 39 118 41 120
rect 49 118 51 120
rect 49 111 51 113
rect 59 111 61 113
rect 76 104 78 106
rect 115 107 117 109
rect 125 110 127 112
rect 135 118 137 120
rect 145 118 147 120
rect 145 111 147 113
rect 155 111 157 113
rect 172 104 174 106
rect 194 113 196 115
rect 204 113 206 115
rect 214 111 216 113
rect 259 107 261 109
rect 269 110 271 112
rect 279 118 281 120
rect 289 118 291 120
rect 289 111 291 113
rect 299 111 301 113
rect 316 104 318 106
rect 355 107 357 109
rect 365 110 367 112
rect 375 118 377 120
rect 385 118 387 120
rect 385 111 387 113
rect 395 111 397 113
rect 412 104 414 106
rect 434 113 436 115
rect 444 113 446 115
rect 454 111 456 113
rect 506 110 508 112
rect 516 110 518 112
rect 533 110 535 112
rect 550 110 552 112
rect 19 79 21 81
rect 29 77 31 79
rect 39 77 41 79
rect 61 86 63 88
rect 78 79 80 81
rect 88 79 90 81
rect 88 72 90 74
rect 98 72 100 74
rect 108 80 110 82
rect 118 83 120 85
rect 157 86 159 88
rect 174 79 176 81
rect 184 79 186 81
rect 184 72 186 74
rect 194 72 196 74
rect 204 80 206 82
rect 214 83 216 85
rect 258 79 260 81
rect 268 77 270 79
rect 278 77 280 79
rect 300 86 302 88
rect 317 79 319 81
rect 327 79 329 81
rect 327 72 329 74
rect 337 72 339 74
rect 347 80 349 82
rect 357 83 359 85
rect 396 86 398 88
rect 413 79 415 81
rect 423 79 425 81
rect 423 72 425 74
rect 433 72 435 74
rect 443 80 445 82
rect 453 83 455 85
rect 506 80 508 82
rect 516 80 518 82
rect 533 80 535 82
rect 550 80 552 82
rect 19 -37 21 -35
rect 29 -34 31 -32
rect 39 -26 41 -24
rect 49 -26 51 -24
rect 49 -33 51 -31
rect 59 -33 61 -31
rect 76 -40 78 -38
rect 115 -37 117 -35
rect 125 -34 127 -32
rect 135 -26 137 -24
rect 145 -26 147 -24
rect 145 -33 147 -31
rect 155 -33 157 -31
rect 172 -40 174 -38
rect 194 -31 196 -29
rect 204 -31 206 -29
rect 214 -33 216 -31
rect 259 -37 261 -35
rect 269 -34 271 -32
rect 279 -26 281 -24
rect 289 -26 291 -24
rect 289 -33 291 -31
rect 299 -33 301 -31
rect 316 -40 318 -38
rect 355 -37 357 -35
rect 365 -34 367 -32
rect 375 -26 377 -24
rect 385 -26 387 -24
rect 385 -33 387 -31
rect 395 -33 397 -31
rect 412 -40 414 -38
rect 434 -31 436 -29
rect 444 -31 446 -29
rect 454 -33 456 -31
rect 506 -34 508 -32
rect 516 -34 518 -32
rect 533 -34 535 -32
rect 550 -34 552 -32
rect 19 -65 21 -63
rect 29 -67 31 -65
rect 39 -67 41 -65
rect 61 -58 63 -56
rect 78 -65 80 -63
rect 88 -65 90 -63
rect 88 -72 90 -70
rect 98 -72 100 -70
rect 108 -64 110 -62
rect 118 -61 120 -59
rect 157 -58 159 -56
rect 174 -65 176 -63
rect 184 -65 186 -63
rect 184 -72 186 -70
rect 194 -72 196 -70
rect 204 -64 206 -62
rect 214 -61 216 -59
rect 258 -65 260 -63
rect 268 -67 270 -65
rect 278 -67 280 -65
rect 300 -58 302 -56
rect 317 -65 319 -63
rect 327 -65 329 -63
rect 327 -72 329 -70
rect 337 -72 339 -70
rect 347 -64 349 -62
rect 357 -61 359 -59
rect 396 -58 398 -56
rect 413 -65 415 -63
rect 423 -65 425 -63
rect 423 -72 425 -70
rect 433 -72 435 -70
rect 443 -64 445 -62
rect 453 -61 455 -59
rect 506 -64 508 -62
rect 516 -64 518 -62
rect 533 -64 535 -62
rect 550 -64 552 -62
<< ndifct1 >>
rect 86 233 88 235
rect 24 223 26 225
rect 24 216 26 218
rect 57 223 59 225
rect 109 233 111 235
rect 98 223 100 225
rect 57 216 59 218
rect 118 221 120 223
rect 148 223 150 225
rect 148 216 150 218
rect 194 223 196 225
rect 268 224 270 226
rect 194 216 196 218
rect 297 216 299 218
rect 378 224 380 226
rect 412 223 414 225
rect 464 223 466 225
rect 506 223 508 225
rect 550 223 552 225
rect 9 111 11 113
rect 87 111 89 113
rect 105 111 107 113
rect 183 111 185 113
rect 224 118 226 120
rect 224 111 226 113
rect 249 111 251 113
rect 327 111 329 113
rect 345 111 347 113
rect 423 111 425 113
rect 464 118 466 120
rect 464 111 466 113
rect 560 110 562 112
rect 9 79 11 81
rect 9 72 11 74
rect 50 79 52 81
rect 128 79 130 81
rect 146 79 148 81
rect 224 79 226 81
rect 248 79 250 81
rect 248 72 250 74
rect 289 79 291 81
rect 367 79 369 81
rect 385 79 387 81
rect 463 79 465 81
rect 560 80 562 82
rect 9 -33 11 -31
rect 87 -33 89 -31
rect 105 -33 107 -31
rect 183 -33 185 -31
rect 224 -26 226 -24
rect 224 -33 226 -31
rect 249 -33 251 -31
rect 327 -33 329 -31
rect 345 -33 347 -31
rect 423 -33 425 -31
rect 464 -26 466 -24
rect 464 -33 466 -31
rect 560 -34 562 -32
rect 9 -65 11 -63
rect 9 -72 11 -70
rect 50 -65 52 -63
rect 128 -65 130 -63
rect 146 -65 148 -63
rect 224 -65 226 -63
rect 248 -65 250 -63
rect 248 -72 250 -70
rect 289 -65 291 -63
rect 367 -65 369 -63
rect 385 -65 387 -63
rect 463 -65 465 -63
rect 560 -64 562 -62
<< ntiect1 >>
rect 127 173 129 175
rect 215 173 217 175
rect 325 173 327 175
rect 507 161 509 163
rect 507 29 509 31
rect 507 17 509 19
rect 507 -115 509 -113
<< ptiect1 >>
rect 119 233 121 235
rect 127 233 129 235
rect 286 233 288 235
rect 197 101 199 103
rect 437 101 439 103
rect 36 89 38 91
rect 275 89 277 91
rect 197 -43 199 -41
rect 437 -43 439 -41
rect 36 -55 38 -53
rect 275 -55 277 -53
<< pdifct0 >>
rect 14 183 16 185
rect 14 176 16 178
rect 47 183 49 185
rect 47 176 49 178
rect 88 184 90 186
rect 88 176 90 178
rect 158 183 160 185
rect 158 176 160 178
rect 184 183 186 185
rect 184 176 186 178
rect 214 198 216 200
rect 224 184 226 186
rect 241 190 243 192
rect 258 184 260 186
rect 287 183 289 185
rect 287 176 289 178
rect 297 183 299 185
rect 324 198 326 200
rect 392 198 394 200
rect 307 183 309 185
rect 334 184 336 186
rect 351 190 353 192
rect 368 184 370 186
rect 392 191 394 193
rect 307 176 309 178
rect 402 183 404 185
rect 402 176 404 178
rect 444 198 446 200
rect 444 191 446 193
rect 422 183 424 185
rect 422 176 424 178
rect 454 183 456 185
rect 454 176 456 178
rect 486 198 488 200
rect 486 191 488 193
rect 474 183 476 185
rect 474 176 476 178
rect 496 183 498 185
rect 496 176 498 178
rect 530 198 532 200
rect 530 191 532 193
rect 516 183 518 185
rect 516 176 518 178
rect 540 183 542 185
rect 540 176 542 178
rect 560 183 562 185
rect 560 176 562 178
rect 20 158 22 160
rect 32 139 34 141
rect 55 158 57 160
rect 55 151 57 153
rect 67 150 69 152
rect 67 143 69 145
rect 77 158 79 160
rect 77 151 79 153
rect 116 158 118 160
rect 128 139 130 141
rect 151 158 153 160
rect 151 151 153 153
rect 163 150 165 152
rect 163 143 165 145
rect 173 158 175 160
rect 173 151 175 153
rect 194 152 196 154
rect 260 158 262 160
rect 272 139 274 141
rect 295 158 297 160
rect 295 151 297 153
rect 307 150 309 152
rect 307 143 309 145
rect 317 158 319 160
rect 317 151 319 153
rect 356 158 358 160
rect 368 139 370 141
rect 391 158 393 160
rect 391 151 393 153
rect 403 150 405 152
rect 403 143 405 145
rect 413 158 415 160
rect 413 151 415 153
rect 434 152 436 154
rect 516 150 518 152
rect 533 144 535 146
rect 550 150 552 152
rect 506 136 508 138
rect 39 38 41 40
rect 60 39 62 41
rect 60 32 62 34
rect 70 47 72 49
rect 70 40 72 42
rect 82 39 84 41
rect 82 32 84 34
rect 105 51 107 53
rect 117 32 119 34
rect 156 39 158 41
rect 156 32 158 34
rect 166 47 168 49
rect 166 40 168 42
rect 178 39 180 41
rect 178 32 180 34
rect 201 51 203 53
rect 213 32 215 34
rect 278 38 280 40
rect 299 39 301 41
rect 299 32 301 34
rect 309 47 311 49
rect 309 40 311 42
rect 321 39 323 41
rect 321 32 323 34
rect 344 51 346 53
rect 356 32 358 34
rect 395 39 397 41
rect 395 32 397 34
rect 405 47 407 49
rect 405 40 407 42
rect 417 39 419 41
rect 417 32 419 34
rect 440 51 442 53
rect 452 32 454 34
rect 506 54 508 56
rect 516 40 518 42
rect 533 46 535 48
rect 550 40 552 42
rect 20 14 22 16
rect 32 -5 34 -3
rect 55 14 57 16
rect 55 7 57 9
rect 67 6 69 8
rect 67 -1 69 1
rect 77 14 79 16
rect 77 7 79 9
rect 116 14 118 16
rect 128 -5 130 -3
rect 151 14 153 16
rect 151 7 153 9
rect 163 6 165 8
rect 163 -1 165 1
rect 173 14 175 16
rect 173 7 175 9
rect 194 8 196 10
rect 260 14 262 16
rect 272 -5 274 -3
rect 295 14 297 16
rect 295 7 297 9
rect 307 6 309 8
rect 307 -1 309 1
rect 317 14 319 16
rect 317 7 319 9
rect 356 14 358 16
rect 368 -5 370 -3
rect 391 14 393 16
rect 391 7 393 9
rect 403 6 405 8
rect 403 -1 405 1
rect 413 14 415 16
rect 413 7 415 9
rect 434 8 436 10
rect 516 6 518 8
rect 533 0 535 2
rect 550 6 552 8
rect 506 -8 508 -6
rect 39 -106 41 -104
rect 60 -105 62 -103
rect 60 -112 62 -110
rect 70 -97 72 -95
rect 70 -104 72 -102
rect 82 -105 84 -103
rect 82 -112 84 -110
rect 105 -93 107 -91
rect 117 -112 119 -110
rect 156 -105 158 -103
rect 156 -112 158 -110
rect 166 -97 168 -95
rect 166 -104 168 -102
rect 178 -105 180 -103
rect 178 -112 180 -110
rect 201 -93 203 -91
rect 213 -112 215 -110
rect 278 -106 280 -104
rect 299 -105 301 -103
rect 299 -112 301 -110
rect 309 -97 311 -95
rect 309 -104 311 -102
rect 321 -105 323 -103
rect 321 -112 323 -110
rect 344 -93 346 -91
rect 356 -112 358 -110
rect 395 -105 397 -103
rect 395 -112 397 -110
rect 405 -97 407 -95
rect 405 -104 407 -102
rect 417 -105 419 -103
rect 417 -112 419 -110
rect 440 -93 442 -91
rect 452 -112 454 -110
rect 506 -90 508 -88
rect 516 -104 518 -102
rect 533 -98 535 -96
rect 550 -104 552 -102
<< pdifct1 >>
rect 24 197 26 199
rect 24 190 26 192
rect 57 197 59 199
rect 148 197 150 199
rect 57 190 59 192
rect 148 190 150 192
rect 119 183 121 185
rect 194 197 196 199
rect 194 190 196 192
rect 268 190 270 192
rect 297 190 299 192
rect 378 190 380 192
rect 412 190 414 192
rect 412 183 414 185
rect 464 190 466 192
rect 464 183 466 185
rect 506 190 508 192
rect 506 183 508 185
rect 550 190 552 192
rect 550 183 552 185
rect 9 146 11 148
rect 9 139 11 141
rect 87 143 89 145
rect 87 136 89 138
rect 105 146 107 148
rect 105 139 107 141
rect 183 143 185 145
rect 183 136 185 138
rect 213 161 215 163
rect 224 152 226 154
rect 224 145 226 147
rect 249 146 251 148
rect 249 139 251 141
rect 327 143 329 145
rect 327 136 329 138
rect 345 146 347 148
rect 345 139 347 141
rect 423 143 425 145
rect 423 136 425 138
rect 453 161 455 163
rect 464 152 466 154
rect 464 145 466 147
rect 560 144 562 146
rect 9 45 11 47
rect 9 38 11 40
rect 20 29 22 31
rect 50 54 52 56
rect 50 47 52 49
rect 128 51 130 53
rect 128 44 130 46
rect 146 54 148 56
rect 146 47 148 49
rect 224 51 226 53
rect 224 44 226 46
rect 248 45 250 47
rect 248 38 250 40
rect 259 29 261 31
rect 289 54 291 56
rect 289 47 291 49
rect 367 51 369 53
rect 367 44 369 46
rect 385 54 387 56
rect 385 47 387 49
rect 463 51 465 53
rect 463 44 465 46
rect 560 46 562 48
rect 9 2 11 4
rect 9 -5 11 -3
rect 87 -1 89 1
rect 87 -8 89 -6
rect 105 2 107 4
rect 105 -5 107 -3
rect 183 -1 185 1
rect 183 -8 185 -6
rect 213 17 215 19
rect 224 8 226 10
rect 224 1 226 3
rect 249 2 251 4
rect 249 -5 251 -3
rect 327 -1 329 1
rect 327 -8 329 -6
rect 345 2 347 4
rect 345 -5 347 -3
rect 423 -1 425 1
rect 423 -8 425 -6
rect 453 17 455 19
rect 464 8 466 10
rect 464 1 466 3
rect 560 0 562 2
rect 9 -99 11 -97
rect 9 -106 11 -104
rect 20 -115 22 -113
rect 50 -90 52 -88
rect 50 -97 52 -95
rect 128 -93 130 -91
rect 128 -100 130 -98
rect 146 -90 148 -88
rect 146 -97 148 -95
rect 224 -93 226 -91
rect 224 -100 226 -98
rect 248 -99 250 -97
rect 248 -106 250 -104
rect 259 -115 261 -113
rect 289 -90 291 -88
rect 289 -97 291 -95
rect 367 -93 369 -91
rect 367 -100 369 -98
rect 385 -90 387 -88
rect 385 -97 387 -95
rect 463 -93 465 -91
rect 463 -100 465 -98
rect 560 -98 562 -96
<< alu0 >>
rect 13 226 17 232
rect 13 224 14 226
rect 16 224 17 226
rect 13 219 17 224
rect 13 217 14 219
rect 16 217 17 219
rect 13 215 17 217
rect 23 214 24 227
rect 46 226 50 232
rect 46 224 47 226
rect 49 224 50 226
rect 46 219 50 224
rect 46 217 47 219
rect 49 217 50 219
rect 46 215 50 217
rect 56 214 57 227
rect 23 195 24 201
rect 56 195 57 201
rect 127 223 131 232
rect 127 221 128 223
rect 130 221 131 223
rect 127 219 131 221
rect 99 213 105 214
rect 110 209 114 211
rect 110 207 111 209
rect 113 207 114 209
rect 110 202 114 207
rect 112 198 114 202
rect 87 186 91 188
rect 12 185 18 186
rect 12 183 14 185
rect 16 183 18 185
rect 12 178 18 183
rect 12 176 14 178
rect 16 176 18 178
rect 45 185 51 186
rect 45 183 47 185
rect 49 183 51 185
rect 45 178 51 183
rect 45 176 47 178
rect 49 176 51 178
rect 87 184 88 186
rect 90 184 91 186
rect 87 178 91 184
rect 150 214 151 227
rect 157 226 161 232
rect 157 224 158 226
rect 160 224 161 226
rect 157 219 161 224
rect 157 217 158 219
rect 160 217 161 219
rect 157 215 161 217
rect 183 226 187 232
rect 183 224 184 226
rect 186 224 187 226
rect 183 219 187 224
rect 183 217 184 219
rect 186 217 187 219
rect 183 215 187 217
rect 193 214 194 227
rect 150 195 151 201
rect 193 195 194 201
rect 212 226 218 227
rect 212 224 214 226
rect 216 224 218 226
rect 212 223 218 224
rect 222 226 228 232
rect 222 224 224 226
rect 226 224 228 226
rect 222 223 228 224
rect 239 226 254 227
rect 239 224 241 226
rect 243 224 254 226
rect 239 223 254 224
rect 212 201 216 223
rect 250 219 254 223
rect 257 226 261 232
rect 257 224 258 226
rect 260 224 261 226
rect 257 222 261 224
rect 236 217 247 219
rect 236 215 244 217
rect 246 215 247 217
rect 250 217 265 219
rect 250 215 262 217
rect 264 215 265 217
rect 236 213 247 215
rect 236 201 240 213
rect 212 200 237 201
rect 212 198 214 200
rect 216 199 237 200
rect 239 199 240 201
rect 216 198 240 199
rect 261 201 265 215
rect 212 197 240 198
rect 252 197 265 201
rect 286 222 290 232
rect 306 229 310 232
rect 306 227 307 229
rect 309 227 310 229
rect 306 225 310 227
rect 322 226 328 227
rect 286 220 287 222
rect 289 220 290 222
rect 286 218 290 220
rect 322 224 324 226
rect 326 224 328 226
rect 322 223 328 224
rect 332 226 338 232
rect 332 224 334 226
rect 336 224 338 226
rect 332 223 338 224
rect 349 226 364 227
rect 349 224 351 226
rect 353 224 364 226
rect 349 223 364 224
rect 252 194 256 197
rect 322 201 326 223
rect 360 219 364 223
rect 367 226 371 232
rect 401 227 405 232
rect 421 227 425 232
rect 453 227 457 232
rect 473 227 477 232
rect 495 227 499 232
rect 515 227 519 232
rect 539 227 543 232
rect 559 227 563 232
rect 367 224 368 226
rect 370 224 371 226
rect 367 222 371 224
rect 346 217 357 219
rect 346 215 354 217
rect 356 215 357 217
rect 360 217 375 219
rect 360 215 372 217
rect 374 215 375 217
rect 346 213 357 215
rect 346 201 350 213
rect 322 200 347 201
rect 322 198 324 200
rect 326 199 347 200
rect 349 199 350 201
rect 326 198 350 199
rect 371 201 375 215
rect 322 197 350 198
rect 362 197 375 201
rect 362 194 366 197
rect 239 192 256 194
rect 239 190 241 192
rect 243 190 256 192
rect 239 189 245 190
rect 156 185 162 186
rect 156 183 158 185
rect 160 183 162 185
rect 87 176 88 178
rect 90 176 91 178
rect 156 178 162 183
rect 156 176 158 178
rect 160 176 162 178
rect 182 185 188 186
rect 182 183 184 185
rect 186 183 188 185
rect 182 178 188 183
rect 222 186 228 187
rect 222 184 224 186
rect 226 184 228 186
rect 182 176 184 178
rect 186 176 188 178
rect 222 176 228 184
rect 256 186 262 187
rect 256 184 258 186
rect 260 184 262 186
rect 256 176 262 184
rect 285 185 291 186
rect 285 183 287 185
rect 289 183 291 185
rect 285 178 291 183
rect 296 185 300 190
rect 349 192 366 194
rect 349 190 351 192
rect 353 190 366 192
rect 349 189 355 190
rect 390 226 396 227
rect 390 224 392 226
rect 394 224 396 226
rect 390 219 396 224
rect 401 225 402 227
rect 404 225 405 227
rect 401 223 405 225
rect 390 217 392 219
rect 394 218 396 219
rect 394 217 411 218
rect 390 214 411 217
rect 390 202 394 214
rect 407 210 411 214
rect 407 208 408 210
rect 410 208 411 210
rect 407 206 411 208
rect 421 225 422 227
rect 424 225 425 227
rect 421 219 425 225
rect 421 217 422 219
rect 424 217 425 219
rect 421 215 425 217
rect 442 226 448 227
rect 442 224 444 226
rect 446 224 448 226
rect 442 219 448 224
rect 453 225 454 227
rect 456 225 457 227
rect 453 223 457 225
rect 442 217 444 219
rect 446 218 448 219
rect 446 217 463 218
rect 442 214 463 217
rect 390 200 395 202
rect 390 198 392 200
rect 394 198 395 200
rect 390 193 395 198
rect 390 191 392 193
rect 394 191 395 193
rect 390 189 395 191
rect 442 202 446 214
rect 459 210 463 214
rect 459 208 460 210
rect 462 208 463 210
rect 459 206 463 208
rect 473 225 474 227
rect 476 225 477 227
rect 473 219 477 225
rect 473 217 474 219
rect 476 217 477 219
rect 473 215 477 217
rect 484 226 490 227
rect 484 224 486 226
rect 488 224 490 226
rect 484 219 490 224
rect 495 225 496 227
rect 498 225 499 227
rect 495 223 499 225
rect 484 217 486 219
rect 488 218 490 219
rect 488 217 505 218
rect 484 214 505 217
rect 442 200 447 202
rect 442 198 444 200
rect 446 198 447 200
rect 442 193 447 198
rect 442 191 444 193
rect 446 191 447 193
rect 296 183 297 185
rect 299 183 300 185
rect 296 181 300 183
rect 305 185 311 186
rect 305 183 307 185
rect 309 183 311 185
rect 285 176 287 178
rect 289 176 291 178
rect 305 178 311 183
rect 332 186 338 187
rect 332 184 334 186
rect 336 184 338 186
rect 305 176 307 178
rect 309 176 311 178
rect 332 176 338 184
rect 366 186 372 187
rect 366 184 368 186
rect 370 184 372 186
rect 366 176 372 184
rect 400 185 406 186
rect 400 183 402 185
rect 404 183 406 185
rect 400 178 406 183
rect 442 189 447 191
rect 484 202 488 214
rect 501 210 505 214
rect 501 208 502 210
rect 504 208 505 210
rect 501 206 505 208
rect 515 225 516 227
rect 518 225 519 227
rect 515 219 519 225
rect 515 217 516 219
rect 518 217 519 219
rect 515 215 519 217
rect 528 226 534 227
rect 528 224 530 226
rect 532 224 534 226
rect 528 219 534 224
rect 539 225 540 227
rect 542 225 543 227
rect 539 223 543 225
rect 528 217 530 219
rect 532 218 534 219
rect 532 217 549 218
rect 528 214 549 217
rect 484 200 489 202
rect 484 198 486 200
rect 488 198 489 200
rect 484 193 489 198
rect 484 191 486 193
rect 488 191 489 193
rect 420 185 426 186
rect 420 183 422 185
rect 424 183 426 185
rect 400 176 402 178
rect 404 176 406 178
rect 420 178 426 183
rect 420 176 422 178
rect 424 176 426 178
rect 452 185 458 186
rect 452 183 454 185
rect 456 183 458 185
rect 452 178 458 183
rect 484 189 489 191
rect 528 202 532 214
rect 545 210 549 214
rect 545 208 546 210
rect 548 208 549 210
rect 545 206 549 208
rect 559 225 560 227
rect 562 225 563 227
rect 559 219 563 225
rect 559 217 560 219
rect 562 217 563 219
rect 559 215 563 217
rect 528 200 533 202
rect 528 198 530 200
rect 532 198 533 200
rect 528 193 533 198
rect 528 191 530 193
rect 532 191 533 193
rect 472 185 478 186
rect 472 183 474 185
rect 476 183 478 185
rect 452 176 454 178
rect 456 176 458 178
rect 472 178 478 183
rect 472 176 474 178
rect 476 176 478 178
rect 494 185 500 186
rect 494 183 496 185
rect 498 183 500 185
rect 494 178 500 183
rect 528 189 533 191
rect 514 185 520 186
rect 514 183 516 185
rect 518 183 520 185
rect 494 176 496 178
rect 498 176 500 178
rect 514 178 520 183
rect 514 176 516 178
rect 518 176 520 178
rect 538 185 544 186
rect 538 183 540 185
rect 542 183 544 185
rect 538 178 544 183
rect 558 185 564 186
rect 558 183 560 185
rect 562 183 564 185
rect 538 176 540 178
rect 542 176 544 178
rect 558 178 564 183
rect 558 176 560 178
rect 562 176 564 178
rect 18 158 20 160
rect 22 158 24 160
rect 18 157 24 158
rect 53 158 55 160
rect 57 158 59 160
rect 53 153 59 158
rect 75 158 77 160
rect 79 158 81 160
rect 53 151 55 153
rect 57 151 59 153
rect 53 150 59 151
rect 66 152 70 154
rect 66 150 67 152
rect 69 150 70 152
rect 75 153 81 158
rect 114 158 116 160
rect 118 158 120 160
rect 114 157 120 158
rect 149 158 151 160
rect 153 158 155 160
rect 75 151 77 153
rect 79 151 81 153
rect 75 150 81 151
rect 149 153 155 158
rect 171 158 173 160
rect 175 158 177 160
rect 149 151 151 153
rect 153 151 155 153
rect 149 150 155 151
rect 162 152 166 154
rect 162 150 163 152
rect 165 150 166 152
rect 171 153 177 158
rect 258 158 260 160
rect 262 158 264 160
rect 258 157 264 158
rect 293 158 295 160
rect 297 158 299 160
rect 171 151 173 153
rect 175 151 177 153
rect 192 154 212 155
rect 192 152 194 154
rect 196 152 212 154
rect 192 151 212 152
rect 171 150 177 151
rect 23 146 47 150
rect 66 146 70 150
rect 21 142 27 146
rect 43 145 83 146
rect 43 143 67 145
rect 69 143 83 145
rect 21 132 25 142
rect 31 141 35 143
rect 43 142 83 143
rect 31 139 32 141
rect 34 139 35 141
rect 31 138 35 139
rect 21 130 22 132
rect 24 130 25 132
rect 21 128 25 130
rect 28 134 35 138
rect 28 123 32 134
rect 71 129 75 134
rect 71 127 72 129
rect 74 127 75 129
rect 14 122 32 123
rect 71 125 75 127
rect 79 131 83 142
rect 79 129 85 131
rect 79 127 82 129
rect 84 127 85 129
rect 79 125 85 127
rect 79 122 83 125
rect 14 120 16 122
rect 18 121 32 122
rect 18 120 43 121
rect 14 119 39 120
rect 28 118 39 119
rect 41 118 43 120
rect 28 117 43 118
rect 48 120 52 122
rect 48 118 49 120
rect 51 118 52 120
rect 48 113 52 118
rect 63 118 83 122
rect 63 114 67 118
rect 119 146 143 150
rect 162 146 166 150
rect 117 142 123 146
rect 139 145 179 146
rect 139 143 163 145
rect 165 143 179 145
rect 117 132 121 142
rect 127 141 131 143
rect 139 142 179 143
rect 127 139 128 141
rect 130 139 131 141
rect 127 138 131 139
rect 117 130 118 132
rect 120 130 121 132
rect 117 128 121 130
rect 124 134 131 138
rect 124 123 128 134
rect 167 129 171 134
rect 167 127 168 129
rect 170 127 171 129
rect 110 122 128 123
rect 110 120 112 122
rect 114 121 128 122
rect 114 120 139 121
rect 110 119 135 120
rect 124 118 135 119
rect 137 118 139 120
rect 124 117 139 118
rect 144 120 148 122
rect 144 118 145 120
rect 147 118 148 120
rect 27 112 49 113
rect 18 109 22 111
rect 27 110 29 112
rect 31 111 49 112
rect 51 111 52 113
rect 31 110 52 111
rect 57 113 67 114
rect 57 111 59 113
rect 61 111 67 113
rect 57 110 67 111
rect 144 113 148 118
rect 167 125 171 127
rect 175 131 179 142
rect 208 146 212 151
rect 208 142 220 146
rect 223 143 224 149
rect 175 129 181 131
rect 175 127 178 129
rect 180 127 181 129
rect 175 125 181 127
rect 175 122 179 125
rect 159 118 179 122
rect 159 114 163 118
rect 196 125 197 141
rect 216 129 220 142
rect 216 127 217 129
rect 219 127 220 129
rect 216 121 220 127
rect 293 153 299 158
rect 315 158 317 160
rect 319 158 321 160
rect 293 151 295 153
rect 297 151 299 153
rect 293 150 299 151
rect 306 152 310 154
rect 306 150 307 152
rect 309 150 310 152
rect 315 153 321 158
rect 354 158 356 160
rect 358 158 360 160
rect 354 157 360 158
rect 389 158 391 160
rect 393 158 395 160
rect 315 151 317 153
rect 319 151 321 153
rect 315 150 321 151
rect 389 153 395 158
rect 411 158 413 160
rect 415 158 417 160
rect 389 151 391 153
rect 393 151 395 153
rect 389 150 395 151
rect 402 152 406 154
rect 402 150 403 152
rect 405 150 406 152
rect 411 153 417 158
rect 411 151 413 153
rect 415 151 417 153
rect 432 154 452 155
rect 432 152 434 154
rect 436 152 452 154
rect 432 151 452 152
rect 411 150 417 151
rect 263 146 287 150
rect 306 146 310 150
rect 261 142 267 146
rect 283 145 323 146
rect 283 143 307 145
rect 309 143 323 145
rect 203 117 220 121
rect 123 112 145 113
rect 27 109 52 110
rect 114 109 118 111
rect 123 110 125 112
rect 127 111 145 112
rect 147 111 148 113
rect 127 110 148 111
rect 153 113 163 114
rect 153 111 155 113
rect 157 111 163 113
rect 153 110 163 111
rect 192 115 198 116
rect 192 113 194 115
rect 196 113 198 115
rect 123 109 148 110
rect 18 107 19 109
rect 21 107 22 109
rect 114 107 115 109
rect 117 107 118 109
rect 18 104 22 107
rect 74 106 80 107
rect 74 104 76 106
rect 78 104 80 106
rect 114 104 118 107
rect 170 106 176 107
rect 170 104 172 106
rect 174 104 176 106
rect 192 104 198 113
rect 203 115 207 117
rect 203 113 204 115
rect 206 113 207 115
rect 203 111 207 113
rect 212 113 218 114
rect 212 111 214 113
rect 216 111 218 113
rect 212 104 218 111
rect 261 132 265 142
rect 271 141 275 143
rect 283 142 323 143
rect 271 139 272 141
rect 274 139 275 141
rect 271 138 275 139
rect 261 130 262 132
rect 264 130 265 132
rect 261 128 265 130
rect 268 134 275 138
rect 268 123 272 134
rect 311 129 315 134
rect 311 127 312 129
rect 314 127 315 129
rect 254 122 272 123
rect 311 125 315 127
rect 319 131 323 142
rect 319 129 325 131
rect 319 127 322 129
rect 324 127 325 129
rect 319 125 325 127
rect 319 122 323 125
rect 254 120 256 122
rect 258 121 272 122
rect 258 120 283 121
rect 254 119 279 120
rect 268 118 279 119
rect 281 118 283 120
rect 268 117 283 118
rect 288 120 292 122
rect 288 118 289 120
rect 291 118 292 120
rect 288 113 292 118
rect 303 118 323 122
rect 303 114 307 118
rect 359 146 383 150
rect 402 146 406 150
rect 357 142 363 146
rect 379 145 419 146
rect 379 143 403 145
rect 405 143 419 145
rect 357 132 361 142
rect 367 141 371 143
rect 379 142 419 143
rect 367 139 368 141
rect 370 139 371 141
rect 367 138 371 139
rect 357 130 358 132
rect 360 130 361 132
rect 357 128 361 130
rect 364 134 371 138
rect 364 123 368 134
rect 407 129 411 134
rect 407 127 408 129
rect 410 127 411 129
rect 350 122 368 123
rect 350 120 352 122
rect 354 121 368 122
rect 354 120 379 121
rect 350 119 375 120
rect 364 118 375 119
rect 377 118 379 120
rect 364 117 379 118
rect 384 120 388 122
rect 384 118 385 120
rect 387 118 388 120
rect 267 112 289 113
rect 258 109 262 111
rect 267 110 269 112
rect 271 111 289 112
rect 291 111 292 113
rect 271 110 292 111
rect 297 113 307 114
rect 297 111 299 113
rect 301 111 307 113
rect 297 110 307 111
rect 384 113 388 118
rect 407 125 411 127
rect 415 131 419 142
rect 448 146 452 151
rect 448 142 460 146
rect 463 143 464 149
rect 415 129 421 131
rect 415 127 418 129
rect 420 127 421 129
rect 415 125 421 127
rect 415 122 419 125
rect 399 118 419 122
rect 399 114 403 118
rect 436 125 437 141
rect 456 129 460 142
rect 456 127 457 129
rect 459 127 460 129
rect 456 121 460 127
rect 514 152 520 160
rect 514 150 516 152
rect 518 150 520 152
rect 514 149 520 150
rect 548 152 554 160
rect 548 150 550 152
rect 552 150 554 152
rect 548 149 554 150
rect 531 146 537 147
rect 531 144 533 146
rect 535 144 548 146
rect 531 142 548 144
rect 544 139 548 142
rect 504 138 532 139
rect 504 136 506 138
rect 508 137 532 138
rect 508 136 529 137
rect 504 135 529 136
rect 531 135 532 137
rect 443 117 460 121
rect 363 112 385 113
rect 267 109 292 110
rect 354 109 358 111
rect 363 110 365 112
rect 367 111 385 112
rect 387 111 388 113
rect 367 110 388 111
rect 393 113 403 114
rect 393 111 395 113
rect 397 111 403 113
rect 393 110 403 111
rect 432 115 438 116
rect 432 113 434 115
rect 436 113 438 115
rect 363 109 388 110
rect 258 107 259 109
rect 261 107 262 109
rect 354 107 355 109
rect 357 107 358 109
rect 258 104 262 107
rect 314 106 320 107
rect 314 104 316 106
rect 318 104 320 106
rect 354 104 358 107
rect 410 106 416 107
rect 410 104 412 106
rect 414 104 416 106
rect 432 104 438 113
rect 443 115 447 117
rect 443 113 444 115
rect 446 113 447 115
rect 443 111 447 113
rect 452 113 458 114
rect 452 111 454 113
rect 456 111 458 113
rect 452 104 458 111
rect 504 113 508 135
rect 528 123 532 135
rect 544 135 557 139
rect 528 121 539 123
rect 553 121 557 135
rect 528 119 536 121
rect 538 119 539 121
rect 528 117 539 119
rect 542 119 554 121
rect 556 119 557 121
rect 542 117 557 119
rect 542 113 546 117
rect 504 112 510 113
rect 504 110 506 112
rect 508 110 510 112
rect 504 109 510 110
rect 514 112 520 113
rect 514 110 516 112
rect 518 110 520 112
rect 514 104 520 110
rect 531 112 546 113
rect 531 110 533 112
rect 535 110 546 112
rect 531 109 546 110
rect 549 112 553 114
rect 549 110 550 112
rect 552 110 553 112
rect 549 104 553 110
rect 17 81 23 88
rect 17 79 19 81
rect 21 79 23 81
rect 17 78 23 79
rect 28 79 32 81
rect 28 77 29 79
rect 31 77 32 79
rect 28 75 32 77
rect 37 79 43 88
rect 59 86 61 88
rect 63 86 65 88
rect 59 85 65 86
rect 117 85 121 88
rect 155 86 157 88
rect 159 86 161 88
rect 155 85 161 86
rect 213 85 217 88
rect 117 83 118 85
rect 120 83 121 85
rect 213 83 214 85
rect 216 83 217 85
rect 87 82 112 83
rect 37 77 39 79
rect 41 77 43 79
rect 37 76 43 77
rect 72 81 82 82
rect 72 79 78 81
rect 80 79 82 81
rect 72 78 82 79
rect 87 81 108 82
rect 87 79 88 81
rect 90 80 108 81
rect 110 80 112 82
rect 117 81 121 83
rect 183 82 208 83
rect 90 79 112 80
rect 15 71 32 75
rect 15 65 19 71
rect 15 63 16 65
rect 18 63 19 65
rect 15 50 19 63
rect 38 51 39 67
rect 72 74 76 78
rect 56 70 76 74
rect 56 67 60 70
rect 54 65 60 67
rect 54 63 55 65
rect 57 63 60 65
rect 54 61 60 63
rect 11 43 12 49
rect 15 46 27 50
rect 23 41 27 46
rect 56 50 60 61
rect 64 65 68 67
rect 87 74 91 79
rect 168 81 178 82
rect 168 79 174 81
rect 176 79 178 81
rect 168 78 178 79
rect 183 81 204 82
rect 183 79 184 81
rect 186 80 204 81
rect 206 80 208 82
rect 213 81 217 83
rect 186 79 208 80
rect 87 72 88 74
rect 90 72 91 74
rect 87 70 91 72
rect 96 74 111 75
rect 96 72 98 74
rect 100 73 111 74
rect 100 72 125 73
rect 96 71 121 72
rect 107 70 121 71
rect 123 70 125 72
rect 107 69 125 70
rect 64 63 65 65
rect 67 63 68 65
rect 64 58 68 63
rect 107 58 111 69
rect 104 54 111 58
rect 114 62 118 64
rect 114 60 115 62
rect 117 60 118 62
rect 104 53 108 54
rect 104 51 105 53
rect 107 51 108 53
rect 56 49 96 50
rect 104 49 108 51
rect 114 50 118 60
rect 56 47 70 49
rect 72 47 96 49
rect 56 46 96 47
rect 112 46 118 50
rect 69 42 73 46
rect 92 42 116 46
rect 168 74 172 78
rect 152 70 172 74
rect 183 74 187 79
rect 183 72 184 74
rect 186 72 187 74
rect 183 70 187 72
rect 192 74 207 75
rect 192 72 194 74
rect 196 73 207 74
rect 196 72 221 73
rect 192 71 217 72
rect 203 70 217 71
rect 219 70 221 72
rect 152 67 156 70
rect 150 65 156 67
rect 150 63 151 65
rect 153 63 156 65
rect 150 61 156 63
rect 152 50 156 61
rect 160 65 164 67
rect 203 69 221 70
rect 160 63 161 65
rect 163 63 164 65
rect 160 58 164 63
rect 203 58 207 69
rect 200 54 207 58
rect 210 62 214 64
rect 210 60 211 62
rect 213 60 214 62
rect 200 53 204 54
rect 200 51 201 53
rect 203 51 204 53
rect 152 49 192 50
rect 200 49 204 51
rect 210 50 214 60
rect 256 81 262 88
rect 256 79 258 81
rect 260 79 262 81
rect 256 78 262 79
rect 267 79 271 81
rect 267 77 268 79
rect 270 77 271 79
rect 267 75 271 77
rect 276 79 282 88
rect 298 86 300 88
rect 302 86 304 88
rect 298 85 304 86
rect 356 85 360 88
rect 394 86 396 88
rect 398 86 400 88
rect 394 85 400 86
rect 452 85 456 88
rect 356 83 357 85
rect 359 83 360 85
rect 452 83 453 85
rect 455 83 456 85
rect 326 82 351 83
rect 276 77 278 79
rect 280 77 282 79
rect 276 76 282 77
rect 311 81 321 82
rect 311 79 317 81
rect 319 79 321 81
rect 311 78 321 79
rect 326 81 347 82
rect 326 79 327 81
rect 329 80 347 81
rect 349 80 351 82
rect 356 81 360 83
rect 422 82 447 83
rect 329 79 351 80
rect 254 71 271 75
rect 152 47 166 49
rect 168 47 192 49
rect 152 46 192 47
rect 208 46 214 50
rect 165 42 169 46
rect 188 42 212 46
rect 58 41 64 42
rect 23 40 43 41
rect 23 38 39 40
rect 41 38 43 40
rect 23 37 43 38
rect 58 39 60 41
rect 62 39 64 41
rect 58 34 64 39
rect 69 40 70 42
rect 72 40 73 42
rect 69 38 73 40
rect 80 41 86 42
rect 80 39 82 41
rect 84 39 86 41
rect 58 32 60 34
rect 62 32 64 34
rect 80 34 86 39
rect 154 41 160 42
rect 154 39 156 41
rect 158 39 160 41
rect 80 32 82 34
rect 84 32 86 34
rect 115 34 121 35
rect 115 32 117 34
rect 119 32 121 34
rect 154 34 160 39
rect 165 40 166 42
rect 168 40 169 42
rect 165 38 169 40
rect 176 41 182 42
rect 176 39 178 41
rect 180 39 182 41
rect 154 32 156 34
rect 158 32 160 34
rect 176 34 182 39
rect 254 65 258 71
rect 254 63 255 65
rect 257 63 258 65
rect 254 50 258 63
rect 277 51 278 67
rect 311 74 315 78
rect 295 70 315 74
rect 295 67 299 70
rect 293 65 299 67
rect 293 63 294 65
rect 296 63 299 65
rect 293 61 299 63
rect 250 43 251 49
rect 254 46 266 50
rect 262 41 266 46
rect 295 50 299 61
rect 303 65 307 67
rect 326 74 330 79
rect 407 81 417 82
rect 407 79 413 81
rect 415 79 417 81
rect 407 78 417 79
rect 422 81 443 82
rect 422 79 423 81
rect 425 80 443 81
rect 445 80 447 82
rect 452 81 456 83
rect 425 79 447 80
rect 326 72 327 74
rect 329 72 330 74
rect 326 70 330 72
rect 335 74 350 75
rect 335 72 337 74
rect 339 73 350 74
rect 339 72 364 73
rect 335 71 360 72
rect 346 70 360 71
rect 362 70 364 72
rect 346 69 364 70
rect 303 63 304 65
rect 306 63 307 65
rect 303 58 307 63
rect 346 58 350 69
rect 343 54 350 58
rect 353 62 357 64
rect 353 60 354 62
rect 356 60 357 62
rect 343 53 347 54
rect 343 51 344 53
rect 346 51 347 53
rect 295 49 335 50
rect 343 49 347 51
rect 353 50 357 60
rect 295 47 309 49
rect 311 47 335 49
rect 295 46 335 47
rect 351 46 357 50
rect 308 42 312 46
rect 331 42 355 46
rect 407 74 411 78
rect 391 70 411 74
rect 422 74 426 79
rect 422 72 423 74
rect 425 72 426 74
rect 422 70 426 72
rect 431 74 446 75
rect 431 72 433 74
rect 435 73 446 74
rect 435 72 460 73
rect 431 71 456 72
rect 442 70 456 71
rect 458 70 460 72
rect 391 67 395 70
rect 389 65 395 67
rect 389 63 390 65
rect 392 63 395 65
rect 389 61 395 63
rect 391 50 395 61
rect 399 65 403 67
rect 442 69 460 70
rect 399 63 400 65
rect 402 63 403 65
rect 399 58 403 63
rect 442 58 446 69
rect 439 54 446 58
rect 449 62 453 64
rect 449 60 450 62
rect 452 60 453 62
rect 439 53 443 54
rect 439 51 440 53
rect 442 51 443 53
rect 391 49 431 50
rect 439 49 443 51
rect 449 50 453 60
rect 391 47 405 49
rect 407 47 431 49
rect 391 46 431 47
rect 447 46 453 50
rect 504 82 510 83
rect 504 80 506 82
rect 508 80 510 82
rect 504 79 510 80
rect 514 82 520 88
rect 514 80 516 82
rect 518 80 520 82
rect 514 79 520 80
rect 531 82 546 83
rect 531 80 533 82
rect 535 80 546 82
rect 531 79 546 80
rect 504 57 508 79
rect 542 75 546 79
rect 549 82 553 88
rect 549 80 550 82
rect 552 80 553 82
rect 549 78 553 80
rect 528 73 539 75
rect 528 71 536 73
rect 538 71 539 73
rect 542 73 557 75
rect 542 71 554 73
rect 556 71 557 73
rect 528 69 539 71
rect 528 57 532 69
rect 504 56 529 57
rect 504 54 506 56
rect 508 55 529 56
rect 531 55 532 57
rect 508 54 532 55
rect 553 57 557 71
rect 504 53 532 54
rect 544 53 557 57
rect 544 50 548 53
rect 404 42 408 46
rect 427 42 451 46
rect 297 41 303 42
rect 262 40 282 41
rect 262 38 278 40
rect 280 38 282 40
rect 262 37 282 38
rect 297 39 299 41
rect 301 39 303 41
rect 176 32 178 34
rect 180 32 182 34
rect 211 34 217 35
rect 211 32 213 34
rect 215 32 217 34
rect 297 34 303 39
rect 308 40 309 42
rect 311 40 312 42
rect 308 38 312 40
rect 319 41 325 42
rect 319 39 321 41
rect 323 39 325 41
rect 297 32 299 34
rect 301 32 303 34
rect 319 34 325 39
rect 393 41 399 42
rect 393 39 395 41
rect 397 39 399 41
rect 319 32 321 34
rect 323 32 325 34
rect 354 34 360 35
rect 354 32 356 34
rect 358 32 360 34
rect 393 34 399 39
rect 404 40 405 42
rect 407 40 408 42
rect 404 38 408 40
rect 415 41 421 42
rect 415 39 417 41
rect 419 39 421 41
rect 393 32 395 34
rect 397 32 399 34
rect 415 34 421 39
rect 531 48 548 50
rect 531 46 533 48
rect 535 46 548 48
rect 531 45 537 46
rect 514 42 520 43
rect 514 40 516 42
rect 518 40 520 42
rect 415 32 417 34
rect 419 32 421 34
rect 450 34 456 35
rect 450 32 452 34
rect 454 32 456 34
rect 514 32 520 40
rect 548 42 554 43
rect 548 40 550 42
rect 552 40 554 42
rect 548 32 554 40
rect 18 14 20 16
rect 22 14 24 16
rect 18 13 24 14
rect 53 14 55 16
rect 57 14 59 16
rect 53 9 59 14
rect 75 14 77 16
rect 79 14 81 16
rect 53 7 55 9
rect 57 7 59 9
rect 53 6 59 7
rect 66 8 70 10
rect 66 6 67 8
rect 69 6 70 8
rect 75 9 81 14
rect 114 14 116 16
rect 118 14 120 16
rect 114 13 120 14
rect 149 14 151 16
rect 153 14 155 16
rect 75 7 77 9
rect 79 7 81 9
rect 75 6 81 7
rect 149 9 155 14
rect 171 14 173 16
rect 175 14 177 16
rect 149 7 151 9
rect 153 7 155 9
rect 149 6 155 7
rect 162 8 166 10
rect 162 6 163 8
rect 165 6 166 8
rect 171 9 177 14
rect 258 14 260 16
rect 262 14 264 16
rect 258 13 264 14
rect 293 14 295 16
rect 297 14 299 16
rect 171 7 173 9
rect 175 7 177 9
rect 192 10 212 11
rect 192 8 194 10
rect 196 8 212 10
rect 192 7 212 8
rect 171 6 177 7
rect 23 2 47 6
rect 66 2 70 6
rect 21 -2 27 2
rect 43 1 83 2
rect 43 -1 67 1
rect 69 -1 83 1
rect 21 -12 25 -2
rect 31 -3 35 -1
rect 43 -2 83 -1
rect 31 -5 32 -3
rect 34 -5 35 -3
rect 31 -6 35 -5
rect 21 -14 22 -12
rect 24 -14 25 -12
rect 21 -16 25 -14
rect 28 -10 35 -6
rect 28 -21 32 -10
rect 71 -15 75 -10
rect 71 -17 72 -15
rect 74 -17 75 -15
rect 14 -22 32 -21
rect 71 -19 75 -17
rect 79 -13 83 -2
rect 79 -15 85 -13
rect 79 -17 82 -15
rect 84 -17 85 -15
rect 79 -19 85 -17
rect 79 -22 83 -19
rect 14 -24 16 -22
rect 18 -23 32 -22
rect 18 -24 43 -23
rect 14 -25 39 -24
rect 28 -26 39 -25
rect 41 -26 43 -24
rect 28 -27 43 -26
rect 48 -24 52 -22
rect 48 -26 49 -24
rect 51 -26 52 -24
rect 48 -31 52 -26
rect 63 -26 83 -22
rect 63 -30 67 -26
rect 119 2 143 6
rect 162 2 166 6
rect 117 -2 123 2
rect 139 1 179 2
rect 139 -1 163 1
rect 165 -1 179 1
rect 117 -12 121 -2
rect 127 -3 131 -1
rect 139 -2 179 -1
rect 127 -5 128 -3
rect 130 -5 131 -3
rect 127 -6 131 -5
rect 117 -14 118 -12
rect 120 -14 121 -12
rect 117 -16 121 -14
rect 124 -10 131 -6
rect 124 -21 128 -10
rect 167 -15 171 -10
rect 167 -17 168 -15
rect 170 -17 171 -15
rect 110 -22 128 -21
rect 110 -24 112 -22
rect 114 -23 128 -22
rect 114 -24 139 -23
rect 110 -25 135 -24
rect 124 -26 135 -25
rect 137 -26 139 -24
rect 124 -27 139 -26
rect 144 -24 148 -22
rect 144 -26 145 -24
rect 147 -26 148 -24
rect 27 -32 49 -31
rect 18 -35 22 -33
rect 27 -34 29 -32
rect 31 -33 49 -32
rect 51 -33 52 -31
rect 31 -34 52 -33
rect 57 -31 67 -30
rect 57 -33 59 -31
rect 61 -33 67 -31
rect 57 -34 67 -33
rect 144 -31 148 -26
rect 167 -19 171 -17
rect 175 -13 179 -2
rect 208 2 212 7
rect 208 -2 220 2
rect 223 -1 224 5
rect 175 -15 181 -13
rect 175 -17 178 -15
rect 180 -17 181 -15
rect 175 -19 181 -17
rect 175 -22 179 -19
rect 159 -26 179 -22
rect 159 -30 163 -26
rect 196 -19 197 -3
rect 216 -15 220 -2
rect 216 -17 217 -15
rect 219 -17 220 -15
rect 216 -23 220 -17
rect 293 9 299 14
rect 315 14 317 16
rect 319 14 321 16
rect 293 7 295 9
rect 297 7 299 9
rect 293 6 299 7
rect 306 8 310 10
rect 306 6 307 8
rect 309 6 310 8
rect 315 9 321 14
rect 354 14 356 16
rect 358 14 360 16
rect 354 13 360 14
rect 389 14 391 16
rect 393 14 395 16
rect 315 7 317 9
rect 319 7 321 9
rect 315 6 321 7
rect 389 9 395 14
rect 411 14 413 16
rect 415 14 417 16
rect 389 7 391 9
rect 393 7 395 9
rect 389 6 395 7
rect 402 8 406 10
rect 402 6 403 8
rect 405 6 406 8
rect 411 9 417 14
rect 411 7 413 9
rect 415 7 417 9
rect 432 10 452 11
rect 432 8 434 10
rect 436 8 452 10
rect 432 7 452 8
rect 411 6 417 7
rect 263 2 287 6
rect 306 2 310 6
rect 261 -2 267 2
rect 283 1 323 2
rect 283 -1 307 1
rect 309 -1 323 1
rect 203 -27 220 -23
rect 123 -32 145 -31
rect 27 -35 52 -34
rect 114 -35 118 -33
rect 123 -34 125 -32
rect 127 -33 145 -32
rect 147 -33 148 -31
rect 127 -34 148 -33
rect 153 -31 163 -30
rect 153 -33 155 -31
rect 157 -33 163 -31
rect 153 -34 163 -33
rect 192 -29 198 -28
rect 192 -31 194 -29
rect 196 -31 198 -29
rect 123 -35 148 -34
rect 18 -37 19 -35
rect 21 -37 22 -35
rect 114 -37 115 -35
rect 117 -37 118 -35
rect 18 -40 22 -37
rect 74 -38 80 -37
rect 74 -40 76 -38
rect 78 -40 80 -38
rect 114 -40 118 -37
rect 170 -38 176 -37
rect 170 -40 172 -38
rect 174 -40 176 -38
rect 192 -40 198 -31
rect 203 -29 207 -27
rect 203 -31 204 -29
rect 206 -31 207 -29
rect 203 -33 207 -31
rect 212 -31 218 -30
rect 212 -33 214 -31
rect 216 -33 218 -31
rect 212 -40 218 -33
rect 261 -12 265 -2
rect 271 -3 275 -1
rect 283 -2 323 -1
rect 271 -5 272 -3
rect 274 -5 275 -3
rect 271 -6 275 -5
rect 261 -14 262 -12
rect 264 -14 265 -12
rect 261 -16 265 -14
rect 268 -10 275 -6
rect 268 -21 272 -10
rect 311 -15 315 -10
rect 311 -17 312 -15
rect 314 -17 315 -15
rect 254 -22 272 -21
rect 311 -19 315 -17
rect 319 -13 323 -2
rect 319 -15 325 -13
rect 319 -17 322 -15
rect 324 -17 325 -15
rect 319 -19 325 -17
rect 319 -22 323 -19
rect 254 -24 256 -22
rect 258 -23 272 -22
rect 258 -24 283 -23
rect 254 -25 279 -24
rect 268 -26 279 -25
rect 281 -26 283 -24
rect 268 -27 283 -26
rect 288 -24 292 -22
rect 288 -26 289 -24
rect 291 -26 292 -24
rect 288 -31 292 -26
rect 303 -26 323 -22
rect 303 -30 307 -26
rect 359 2 383 6
rect 402 2 406 6
rect 357 -2 363 2
rect 379 1 419 2
rect 379 -1 403 1
rect 405 -1 419 1
rect 357 -12 361 -2
rect 367 -3 371 -1
rect 379 -2 419 -1
rect 367 -5 368 -3
rect 370 -5 371 -3
rect 367 -6 371 -5
rect 357 -14 358 -12
rect 360 -14 361 -12
rect 357 -16 361 -14
rect 364 -10 371 -6
rect 364 -21 368 -10
rect 407 -15 411 -10
rect 407 -17 408 -15
rect 410 -17 411 -15
rect 350 -22 368 -21
rect 350 -24 352 -22
rect 354 -23 368 -22
rect 354 -24 379 -23
rect 350 -25 375 -24
rect 364 -26 375 -25
rect 377 -26 379 -24
rect 364 -27 379 -26
rect 384 -24 388 -22
rect 384 -26 385 -24
rect 387 -26 388 -24
rect 267 -32 289 -31
rect 258 -35 262 -33
rect 267 -34 269 -32
rect 271 -33 289 -32
rect 291 -33 292 -31
rect 271 -34 292 -33
rect 297 -31 307 -30
rect 297 -33 299 -31
rect 301 -33 307 -31
rect 297 -34 307 -33
rect 384 -31 388 -26
rect 407 -19 411 -17
rect 415 -13 419 -2
rect 448 2 452 7
rect 448 -2 460 2
rect 463 -1 464 5
rect 415 -15 421 -13
rect 415 -17 418 -15
rect 420 -17 421 -15
rect 415 -19 421 -17
rect 415 -22 419 -19
rect 399 -26 419 -22
rect 399 -30 403 -26
rect 436 -19 437 -3
rect 456 -15 460 -2
rect 456 -17 457 -15
rect 459 -17 460 -15
rect 456 -23 460 -17
rect 514 8 520 16
rect 514 6 516 8
rect 518 6 520 8
rect 514 5 520 6
rect 548 8 554 16
rect 548 6 550 8
rect 552 6 554 8
rect 548 5 554 6
rect 531 2 537 3
rect 531 0 533 2
rect 535 0 548 2
rect 531 -2 548 0
rect 544 -5 548 -2
rect 504 -6 532 -5
rect 504 -8 506 -6
rect 508 -7 532 -6
rect 508 -8 529 -7
rect 504 -9 529 -8
rect 531 -9 532 -7
rect 443 -27 460 -23
rect 363 -32 385 -31
rect 267 -35 292 -34
rect 354 -35 358 -33
rect 363 -34 365 -32
rect 367 -33 385 -32
rect 387 -33 388 -31
rect 367 -34 388 -33
rect 393 -31 403 -30
rect 393 -33 395 -31
rect 397 -33 403 -31
rect 393 -34 403 -33
rect 432 -29 438 -28
rect 432 -31 434 -29
rect 436 -31 438 -29
rect 363 -35 388 -34
rect 258 -37 259 -35
rect 261 -37 262 -35
rect 354 -37 355 -35
rect 357 -37 358 -35
rect 258 -40 262 -37
rect 314 -38 320 -37
rect 314 -40 316 -38
rect 318 -40 320 -38
rect 354 -40 358 -37
rect 410 -38 416 -37
rect 410 -40 412 -38
rect 414 -40 416 -38
rect 432 -40 438 -31
rect 443 -29 447 -27
rect 443 -31 444 -29
rect 446 -31 447 -29
rect 443 -33 447 -31
rect 452 -31 458 -30
rect 452 -33 454 -31
rect 456 -33 458 -31
rect 452 -40 458 -33
rect 504 -31 508 -9
rect 528 -21 532 -9
rect 544 -9 557 -5
rect 528 -23 539 -21
rect 553 -23 557 -9
rect 528 -25 536 -23
rect 538 -25 539 -23
rect 528 -27 539 -25
rect 542 -25 554 -23
rect 556 -25 557 -23
rect 542 -27 557 -25
rect 542 -31 546 -27
rect 504 -32 510 -31
rect 504 -34 506 -32
rect 508 -34 510 -32
rect 504 -35 510 -34
rect 514 -32 520 -31
rect 514 -34 516 -32
rect 518 -34 520 -32
rect 514 -40 520 -34
rect 531 -32 546 -31
rect 531 -34 533 -32
rect 535 -34 546 -32
rect 531 -35 546 -34
rect 549 -32 553 -30
rect 549 -34 550 -32
rect 552 -34 553 -32
rect 549 -40 553 -34
rect 17 -63 23 -56
rect 17 -65 19 -63
rect 21 -65 23 -63
rect 17 -66 23 -65
rect 28 -65 32 -63
rect 28 -67 29 -65
rect 31 -67 32 -65
rect 28 -69 32 -67
rect 37 -65 43 -56
rect 59 -58 61 -56
rect 63 -58 65 -56
rect 59 -59 65 -58
rect 117 -59 121 -56
rect 155 -58 157 -56
rect 159 -58 161 -56
rect 155 -59 161 -58
rect 213 -59 217 -56
rect 117 -61 118 -59
rect 120 -61 121 -59
rect 213 -61 214 -59
rect 216 -61 217 -59
rect 87 -62 112 -61
rect 37 -67 39 -65
rect 41 -67 43 -65
rect 37 -68 43 -67
rect 72 -63 82 -62
rect 72 -65 78 -63
rect 80 -65 82 -63
rect 72 -66 82 -65
rect 87 -63 108 -62
rect 87 -65 88 -63
rect 90 -64 108 -63
rect 110 -64 112 -62
rect 117 -63 121 -61
rect 183 -62 208 -61
rect 90 -65 112 -64
rect 15 -73 32 -69
rect 15 -79 19 -73
rect 15 -81 16 -79
rect 18 -81 19 -79
rect 15 -94 19 -81
rect 38 -93 39 -77
rect 72 -70 76 -66
rect 56 -74 76 -70
rect 56 -77 60 -74
rect 54 -79 60 -77
rect 54 -81 55 -79
rect 57 -81 60 -79
rect 54 -83 60 -81
rect 11 -101 12 -95
rect 15 -98 27 -94
rect 23 -103 27 -98
rect 56 -94 60 -83
rect 64 -79 68 -77
rect 87 -70 91 -65
rect 168 -63 178 -62
rect 168 -65 174 -63
rect 176 -65 178 -63
rect 168 -66 178 -65
rect 183 -63 204 -62
rect 183 -65 184 -63
rect 186 -64 204 -63
rect 206 -64 208 -62
rect 213 -63 217 -61
rect 186 -65 208 -64
rect 87 -72 88 -70
rect 90 -72 91 -70
rect 87 -74 91 -72
rect 96 -70 111 -69
rect 96 -72 98 -70
rect 100 -71 111 -70
rect 100 -72 125 -71
rect 96 -73 121 -72
rect 107 -74 121 -73
rect 123 -74 125 -72
rect 107 -75 125 -74
rect 64 -81 65 -79
rect 67 -81 68 -79
rect 64 -86 68 -81
rect 107 -86 111 -75
rect 104 -90 111 -86
rect 114 -82 118 -80
rect 114 -84 115 -82
rect 117 -84 118 -82
rect 104 -91 108 -90
rect 104 -93 105 -91
rect 107 -93 108 -91
rect 56 -95 96 -94
rect 104 -95 108 -93
rect 114 -94 118 -84
rect 56 -97 70 -95
rect 72 -97 96 -95
rect 56 -98 96 -97
rect 112 -98 118 -94
rect 69 -102 73 -98
rect 92 -102 116 -98
rect 168 -70 172 -66
rect 152 -74 172 -70
rect 183 -70 187 -65
rect 183 -72 184 -70
rect 186 -72 187 -70
rect 183 -74 187 -72
rect 192 -70 207 -69
rect 192 -72 194 -70
rect 196 -71 207 -70
rect 196 -72 221 -71
rect 192 -73 217 -72
rect 203 -74 217 -73
rect 219 -74 221 -72
rect 152 -77 156 -74
rect 150 -79 156 -77
rect 150 -81 151 -79
rect 153 -81 156 -79
rect 150 -83 156 -81
rect 152 -94 156 -83
rect 160 -79 164 -77
rect 203 -75 221 -74
rect 160 -81 161 -79
rect 163 -81 164 -79
rect 160 -86 164 -81
rect 203 -86 207 -75
rect 200 -90 207 -86
rect 210 -82 214 -80
rect 210 -84 211 -82
rect 213 -84 214 -82
rect 200 -91 204 -90
rect 200 -93 201 -91
rect 203 -93 204 -91
rect 152 -95 192 -94
rect 200 -95 204 -93
rect 210 -94 214 -84
rect 256 -63 262 -56
rect 256 -65 258 -63
rect 260 -65 262 -63
rect 256 -66 262 -65
rect 267 -65 271 -63
rect 267 -67 268 -65
rect 270 -67 271 -65
rect 267 -69 271 -67
rect 276 -65 282 -56
rect 298 -58 300 -56
rect 302 -58 304 -56
rect 298 -59 304 -58
rect 356 -59 360 -56
rect 394 -58 396 -56
rect 398 -58 400 -56
rect 394 -59 400 -58
rect 452 -59 456 -56
rect 356 -61 357 -59
rect 359 -61 360 -59
rect 452 -61 453 -59
rect 455 -61 456 -59
rect 326 -62 351 -61
rect 276 -67 278 -65
rect 280 -67 282 -65
rect 276 -68 282 -67
rect 311 -63 321 -62
rect 311 -65 317 -63
rect 319 -65 321 -63
rect 311 -66 321 -65
rect 326 -63 347 -62
rect 326 -65 327 -63
rect 329 -64 347 -63
rect 349 -64 351 -62
rect 356 -63 360 -61
rect 422 -62 447 -61
rect 329 -65 351 -64
rect 254 -73 271 -69
rect 152 -97 166 -95
rect 168 -97 192 -95
rect 152 -98 192 -97
rect 208 -98 214 -94
rect 165 -102 169 -98
rect 188 -102 212 -98
rect 58 -103 64 -102
rect 23 -104 43 -103
rect 23 -106 39 -104
rect 41 -106 43 -104
rect 23 -107 43 -106
rect 58 -105 60 -103
rect 62 -105 64 -103
rect 58 -110 64 -105
rect 69 -104 70 -102
rect 72 -104 73 -102
rect 69 -106 73 -104
rect 80 -103 86 -102
rect 80 -105 82 -103
rect 84 -105 86 -103
rect 58 -112 60 -110
rect 62 -112 64 -110
rect 80 -110 86 -105
rect 154 -103 160 -102
rect 154 -105 156 -103
rect 158 -105 160 -103
rect 80 -112 82 -110
rect 84 -112 86 -110
rect 115 -110 121 -109
rect 115 -112 117 -110
rect 119 -112 121 -110
rect 154 -110 160 -105
rect 165 -104 166 -102
rect 168 -104 169 -102
rect 165 -106 169 -104
rect 176 -103 182 -102
rect 176 -105 178 -103
rect 180 -105 182 -103
rect 154 -112 156 -110
rect 158 -112 160 -110
rect 176 -110 182 -105
rect 254 -79 258 -73
rect 254 -81 255 -79
rect 257 -81 258 -79
rect 254 -94 258 -81
rect 277 -93 278 -77
rect 311 -70 315 -66
rect 295 -74 315 -70
rect 295 -77 299 -74
rect 293 -79 299 -77
rect 293 -81 294 -79
rect 296 -81 299 -79
rect 293 -83 299 -81
rect 250 -101 251 -95
rect 254 -98 266 -94
rect 262 -103 266 -98
rect 295 -94 299 -83
rect 303 -79 307 -77
rect 326 -70 330 -65
rect 407 -63 417 -62
rect 407 -65 413 -63
rect 415 -65 417 -63
rect 407 -66 417 -65
rect 422 -63 443 -62
rect 422 -65 423 -63
rect 425 -64 443 -63
rect 445 -64 447 -62
rect 452 -63 456 -61
rect 425 -65 447 -64
rect 326 -72 327 -70
rect 329 -72 330 -70
rect 326 -74 330 -72
rect 335 -70 350 -69
rect 335 -72 337 -70
rect 339 -71 350 -70
rect 339 -72 364 -71
rect 335 -73 360 -72
rect 346 -74 360 -73
rect 362 -74 364 -72
rect 346 -75 364 -74
rect 303 -81 304 -79
rect 306 -81 307 -79
rect 303 -86 307 -81
rect 346 -86 350 -75
rect 343 -90 350 -86
rect 353 -82 357 -80
rect 353 -84 354 -82
rect 356 -84 357 -82
rect 343 -91 347 -90
rect 343 -93 344 -91
rect 346 -93 347 -91
rect 295 -95 335 -94
rect 343 -95 347 -93
rect 353 -94 357 -84
rect 295 -97 309 -95
rect 311 -97 335 -95
rect 295 -98 335 -97
rect 351 -98 357 -94
rect 308 -102 312 -98
rect 331 -102 355 -98
rect 407 -70 411 -66
rect 391 -74 411 -70
rect 422 -70 426 -65
rect 422 -72 423 -70
rect 425 -72 426 -70
rect 422 -74 426 -72
rect 431 -70 446 -69
rect 431 -72 433 -70
rect 435 -71 446 -70
rect 435 -72 460 -71
rect 431 -73 456 -72
rect 442 -74 456 -73
rect 458 -74 460 -72
rect 391 -77 395 -74
rect 389 -79 395 -77
rect 389 -81 390 -79
rect 392 -81 395 -79
rect 389 -83 395 -81
rect 391 -94 395 -83
rect 399 -79 403 -77
rect 442 -75 460 -74
rect 399 -81 400 -79
rect 402 -81 403 -79
rect 399 -86 403 -81
rect 442 -86 446 -75
rect 439 -90 446 -86
rect 449 -82 453 -80
rect 449 -84 450 -82
rect 452 -84 453 -82
rect 439 -91 443 -90
rect 439 -93 440 -91
rect 442 -93 443 -91
rect 391 -95 431 -94
rect 439 -95 443 -93
rect 449 -94 453 -84
rect 391 -97 405 -95
rect 407 -97 431 -95
rect 391 -98 431 -97
rect 447 -98 453 -94
rect 504 -62 510 -61
rect 504 -64 506 -62
rect 508 -64 510 -62
rect 504 -65 510 -64
rect 514 -62 520 -56
rect 514 -64 516 -62
rect 518 -64 520 -62
rect 514 -65 520 -64
rect 531 -62 546 -61
rect 531 -64 533 -62
rect 535 -64 546 -62
rect 531 -65 546 -64
rect 504 -87 508 -65
rect 542 -69 546 -65
rect 549 -62 553 -56
rect 549 -64 550 -62
rect 552 -64 553 -62
rect 549 -66 553 -64
rect 528 -71 539 -69
rect 528 -73 536 -71
rect 538 -73 539 -71
rect 542 -71 557 -69
rect 542 -73 554 -71
rect 556 -73 557 -71
rect 528 -75 539 -73
rect 528 -87 532 -75
rect 504 -88 529 -87
rect 504 -90 506 -88
rect 508 -89 529 -88
rect 531 -89 532 -87
rect 508 -90 532 -89
rect 553 -87 557 -73
rect 504 -91 532 -90
rect 544 -91 557 -87
rect 544 -94 548 -91
rect 404 -102 408 -98
rect 427 -102 451 -98
rect 297 -103 303 -102
rect 262 -104 282 -103
rect 262 -106 278 -104
rect 280 -106 282 -104
rect 262 -107 282 -106
rect 297 -105 299 -103
rect 301 -105 303 -103
rect 176 -112 178 -110
rect 180 -112 182 -110
rect 211 -110 217 -109
rect 211 -112 213 -110
rect 215 -112 217 -110
rect 297 -110 303 -105
rect 308 -104 309 -102
rect 311 -104 312 -102
rect 308 -106 312 -104
rect 319 -103 325 -102
rect 319 -105 321 -103
rect 323 -105 325 -103
rect 297 -112 299 -110
rect 301 -112 303 -110
rect 319 -110 325 -105
rect 393 -103 399 -102
rect 393 -105 395 -103
rect 397 -105 399 -103
rect 319 -112 321 -110
rect 323 -112 325 -110
rect 354 -110 360 -109
rect 354 -112 356 -110
rect 358 -112 360 -110
rect 393 -110 399 -105
rect 404 -104 405 -102
rect 407 -104 408 -102
rect 404 -106 408 -104
rect 415 -103 421 -102
rect 415 -105 417 -103
rect 419 -105 421 -103
rect 393 -112 395 -110
rect 397 -112 399 -110
rect 415 -110 421 -105
rect 531 -96 548 -94
rect 531 -98 533 -96
rect 535 -98 548 -96
rect 531 -99 537 -98
rect 514 -102 520 -101
rect 514 -104 516 -102
rect 518 -104 520 -102
rect 415 -112 417 -110
rect 419 -112 421 -110
rect 450 -110 456 -109
rect 450 -112 452 -110
rect 454 -112 456 -110
rect 514 -112 520 -104
rect 548 -102 554 -101
rect 548 -104 550 -102
rect 552 -104 554 -102
rect 548 -112 554 -104
<< via1 >>
rect 25 203 27 205
rect 88 215 90 217
rect 89 207 91 209
rect 64 190 66 192
rect 117 191 119 193
rect 143 190 145 192
rect 246 199 248 201
rect 197 193 199 195
rect 308 199 310 201
rect 354 199 356 201
rect 97 182 99 184
rect 129 182 131 184
rect 213 182 215 184
rect 423 191 425 193
rect 323 182 325 184
rect 475 191 477 193
rect 517 191 519 193
rect 561 191 563 193
rect 8 151 10 153
rect 56 120 58 122
rect 151 135 153 137
rect 104 120 106 122
rect 96 111 98 113
rect 209 136 211 138
rect 240 130 242 132
rect 248 122 250 124
rect 280 130 282 132
rect 296 120 298 122
rect 376 135 378 137
rect 344 120 346 122
rect 336 111 338 113
rect 449 136 451 138
rect 481 130 483 132
rect 514 120 516 122
rect 9 65 11 67
rect 24 54 26 56
rect 137 79 139 81
rect 129 70 131 72
rect 64 55 66 57
rect 177 70 179 72
rect 225 69 227 71
rect 193 60 195 62
rect 233 60 235 62
rect 263 54 265 56
rect 376 79 378 81
rect 368 70 370 72
rect 308 55 310 57
rect 416 70 418 72
rect 432 60 434 62
rect 517 72 519 74
rect 536 55 538 57
rect 464 41 466 43
rect 56 -24 58 -22
rect 104 -24 106 -22
rect 96 -33 98 -31
rect 209 -8 211 -6
rect 240 -14 242 -12
rect 280 -14 282 -12
rect 296 -24 298 -22
rect 344 -24 346 -22
rect 336 -33 338 -31
rect 449 -8 451 -6
rect 481 -14 483 -12
rect 517 -26 519 -24
rect 536 -9 538 -7
rect 24 -90 26 -88
rect 137 -65 139 -63
rect 129 -74 131 -72
rect 64 -89 66 -87
rect 177 -74 179 -72
rect 193 -84 195 -82
rect 233 -84 235 -82
rect 263 -90 265 -88
rect 376 -65 378 -63
rect 368 -74 370 -72
rect 416 -74 418 -72
rect 432 -84 434 -82
rect 536 -86 538 -84
<< via2 >>
rect 88 215 90 217
rect 89 207 91 209
rect 25 203 27 205
rect 246 199 248 201
rect 197 193 199 195
rect 64 190 66 192
rect 117 191 119 193
rect 143 190 145 192
rect 423 191 425 193
rect 475 191 477 193
rect 517 191 519 193
rect 561 191 563 193
rect 97 182 99 184
rect 129 182 131 184
rect 213 182 215 184
rect 323 182 325 184
rect 8 151 10 153
rect 151 135 153 137
rect 376 135 378 137
rect 248 122 250 124
rect 225 69 227 71
rect 9 65 11 67
rect 514 120 516 122
rect 517 72 519 74
rect 64 55 66 57
rect 308 55 310 57
rect 536 55 538 57
rect 464 41 466 43
rect 536 -9 538 -7
rect 517 -26 519 -24
rect 536 -86 538 -84
rect 64 -89 66 -87
<< via3 >>
rect 8 215 10 217
rect 89 207 91 209
rect 25 203 27 205
rect 246 199 248 201
rect 197 193 199 195
rect 64 190 66 192
rect 117 191 119 193
rect 143 190 145 192
rect 423 191 425 193
rect 475 191 477 193
rect 517 191 519 193
rect 561 191 563 193
rect 97 182 99 184
rect 25 163 27 165
rect 151 163 153 165
rect 8 151 10 153
rect 151 135 153 137
rect 197 135 199 137
rect 117 125 119 127
rect 475 120 477 122
rect 517 72 519 74
rect 89 69 91 71
rect 9 65 11 67
rect 64 55 66 57
rect 143 55 145 57
rect 423 55 425 57
rect 97 41 99 43
rect 25 19 27 21
rect 151 19 153 21
rect 475 -9 477 -7
rect 561 -26 563 -24
rect 517 -86 519 -84
rect 64 -89 66 -87
<< via4 >>
rect 9 65 11 67
rect 246 65 248 67
<< labels >>
rlabel alu1 149 100 149 100 6 vss
rlabel alu1 210 164 210 164 4 vdd
rlabel alu1 210 100 210 100 4 vss
rlabel alu1 153 124 153 124 1 a0
rlabel alu1 161 128 161 128 1 a0
rlabel alu1 218 152 218 152 1 c0
rlabel alu1 226 132 226 132 1 c0
rlabel alu1 389 100 389 100 6 vss
rlabel alu1 389 164 389 164 6 vdd
rlabel alu1 293 164 293 164 6 vdd
rlabel alu1 293 100 293 100 6 vss
rlabel alu1 450 164 450 164 4 vdd
rlabel alu1 450 100 450 100 4 vss
rlabel alu1 297 136 297 136 1 c0
rlabel alu1 393 124 393 124 1 a1
rlabel alu1 401 128 401 128 1 a1
rlabel alu1 458 152 458 152 1 c1
rlabel alu1 466 132 466 132 1 c1
rlabel alu1 53 100 53 100 6 vss
rlabel alu1 325 92 325 92 2 vss
rlabel alu1 325 28 325 28 2 vdd
rlabel alu1 421 28 421 28 2 vdd
rlabel alu1 421 92 421 92 2 vss
rlabel alu1 264 28 264 28 8 vdd
rlabel alu1 264 92 264 92 8 vss
rlabel alu1 417 56 417 56 5 c1
rlabel alu1 321 68 321 68 5 a2
rlabel alu1 313 64 313 64 5 a2
rlabel alu1 256 40 256 40 5 c2
rlabel alu1 248 60 248 60 5 c2
rlabel alu1 86 92 86 92 2 vss
rlabel alu1 86 28 86 28 2 vdd
rlabel alu1 182 28 182 28 2 vdd
rlabel alu1 182 92 182 92 2 vss
rlabel alu1 25 28 25 28 8 vdd
rlabel alu1 25 92 25 92 8 vss
rlabel alu1 178 56 178 56 5 c2
rlabel alu1 82 68 82 68 5 a3
rlabel alu1 74 64 74 64 5 a3
rlabel alu1 17 40 17 40 5 c3
rlabel alu1 9 60 9 60 5 c3
rlabel alu1 153 136 153 136 1 b0i
rlabel alu1 53 164 53 164 6 vdd
rlabel alu1 149 164 149 164 6 vdd
rlabel alu1 26 208 26 208 1 b0i
rlabel alu1 18 192 18 192 1 b0i
rlabel polyct1 18 208 18 208 1 b0
rlabel alu1 10 200 10 200 1 b0
rlabel alu1 18 172 18 172 2 vdd
rlabel alu1 18 236 18 236 2 vss
rlabel alu1 51 236 51 236 2 vss
rlabel alu1 51 172 51 172 2 vdd
rlabel alu1 43 200 43 200 1 b3
rlabel polyct1 51 208 51 208 1 b3
rlabel alu1 51 192 51 192 1 b3i
rlabel alu1 59 208 59 208 1 b3i
rlabel via3 66 56 66 56 1 b3i
rlabel alu1 82 56 82 56 1 b3i
rlabel alu1 106 236 106 236 2 vss
rlabel alu1 106 172 106 172 2 vdd
rlabel alu1 321 56 321 56 1 b2i
rlabel alu1 156 172 156 172 8 vdd
rlabel alu1 156 236 156 236 8 vss
rlabel alu1 164 200 164 200 1 b2
rlabel polyct1 156 208 156 208 1 b2
rlabel alu1 156 192 156 192 1 b2i
rlabel alu1 148 208 148 208 1 b2i
rlabel alu1 188 172 188 172 2 vdd
rlabel alu1 188 236 188 236 2 vss
rlabel alu1 180 200 180 200 1 b1
rlabel polyct1 188 208 188 208 1 b1
rlabel alu1 196 208 196 208 1 b1i
rlabel alu1 188 192 188 192 1 b1i
rlabel alu1 393 136 393 136 1 b1i
rlabel alu1 242 236 242 236 2 vss
rlabel alu1 242 172 242 172 2 vdd
rlabel alu1 270 208 270 208 1 gt
rlabel alu1 262 192 262 192 1 gt
rlabel alu1 246 204 246 204 1 c3
rlabel alu1 254 208 254 208 1 c3
rlabel alu1 222 216 222 216 1 vss
rlabel alu1 230 212 230 212 1 vss
rlabel alu1 352 236 352 236 2 vss
rlabel alu1 352 172 352 172 2 vdd
rlabel alu1 332 216 332 216 1 vss
rlabel alu1 340 212 340 212 1 vss
rlabel alu1 297 172 297 172 2 vdd
rlabel alu1 297 236 297 236 2 vss
rlabel alu1 380 208 380 208 1 lt
rlabel alu1 372 192 372 192 1 lt
rlabel alu1 57 136 57 136 1 c
rlabel alu1 9 128 9 128 1 d0
rlabel alu1 17 152 17 152 1 d0
rlabel alu1 90 220 90 220 1 d0
rlabel alu1 98 216 98 216 1 d0
rlabel alu1 106 216 106 216 1 d0
rlabel alu1 257 152 257 152 1 d1
rlabel alu1 122 200 122 200 1 d1
rlabel alu1 98 208 98 208 1 d3
rlabel alu1 224 39 224 39 1 d3
rlabel alu1 227 48 227 48 1 d3
rlabel alu1 98 188 98 188 1 d2
rlabel alu1 106 200 106 200 1 d2
rlabel alu1 465 64 465 64 1 d2
rlabel alu1 463 39 463 39 1 d2
rlabel alu1 130 196 130 196 1 eq
rlabel alu1 119 216 119 216 1 eq
rlabel alu1 222 192 222 192 1 eq
rlabel alu1 149 -44 149 -44 6 vss
rlabel alu1 65 -8 65 -8 1 cin
rlabel alu1 57 -8 57 -8 1 cin
rlabel alu1 49 -8 49 -8 1 cin
rlabel alu1 41 -12 41 -12 1 cin
rlabel alu1 210 20 210 20 4 vdd
rlabel alu1 210 -44 210 -44 4 vss
rlabel alu1 9 -16 9 -16 1 s0
rlabel alu1 17 8 17 8 1 s0
rlabel alu1 389 -44 389 -44 6 vss
rlabel alu1 389 20 389 20 6 vdd
rlabel alu1 293 20 293 20 6 vdd
rlabel alu1 293 -44 293 -44 6 vss
rlabel alu1 450 20 450 20 4 vdd
rlabel alu1 450 -44 450 -44 4 vss
rlabel alu1 249 -16 249 -16 1 s1
rlabel alu1 257 8 257 8 1 s1
rlabel pmos 73 -8 73 -8 1 cin
rlabel alu1 53 -44 53 -44 6 vss
rlabel alu1 325 -52 325 -52 2 vss
rlabel alu1 325 -116 325 -116 2 vdd
rlabel alu1 421 -116 421 -116 2 vdd
rlabel alu1 421 -52 421 -52 2 vss
rlabel alu1 264 -116 264 -116 8 vdd
rlabel alu1 264 -52 264 -52 8 vss
rlabel alu1 465 -80 465 -80 5 s2
rlabel alu1 457 -104 457 -104 5 s2
rlabel alu1 86 -52 86 -52 2 vss
rlabel alu1 86 -116 86 -116 2 vdd
rlabel alu1 182 -116 182 -116 2 vdd
rlabel alu1 182 -52 182 -52 2 vss
rlabel alu1 25 -116 25 -116 8 vdd
rlabel alu1 25 -52 25 -52 8 vss
rlabel alu1 226 -80 226 -80 5 s3
rlabel alu1 218 -104 218 -104 5 s3
rlabel alu1 53 20 53 20 6 vdd
rlabel alu1 149 20 149 20 6 vdd
rlabel alu1 153 -8 153 -8 1 n0
rlabel alu1 153 -20 153 -20 1 m0
rlabel alu1 218 8 218 8 1 cs0
rlabel alu1 226 -12 226 -12 1 cs0
rlabel alu1 297 -8 297 -8 1 cs0
rlabel alu1 393 -8 393 -8 1 n1
rlabel alu1 393 -20 393 -20 1 m1
rlabel alu1 466 -12 466 -12 1 cs1
rlabel alu1 417 -88 417 -88 1 cs1
rlabel alu1 321 -76 321 -76 1 m2
rlabel alu1 321 -88 321 -88 1 n2
rlabel alu1 248 -84 248 -84 1 cs2
rlabel alu1 178 -88 178 -88 1 cs2
rlabel alu1 82 -88 82 -88 1 n3
rlabel alu1 82 -76 82 -76 1 m3
rlabel alu1 17 -104 17 -104 1 cs3
rlabel alu1 9 -84 9 -84 1 cs3
rlabel alu1 408 236 408 236 2 vss
rlabel alu1 408 172 408 172 2 vdd
rlabel alu1 403 200 403 200 1 p0
rlabel alu1 416 192 416 192 1 q0
rlabel alu1 424 204 424 204 1 q0
rlabel alu1 460 236 460 236 2 vss
rlabel alu1 460 172 460 172 2 vdd
rlabel alu1 455 200 455 200 1 p1
rlabel alu1 476 204 476 204 1 q1
rlabel alu1 468 192 468 192 1 q1
rlabel alu1 502 172 502 172 2 vdd
rlabel alu1 502 236 502 236 2 vss
rlabel alu1 498 200 498 200 1 p2
rlabel alu1 518 204 518 204 1 q2
rlabel alu1 510 192 510 192 1 q2
rlabel alu1 546 236 546 236 2 vss
rlabel alu1 546 172 546 172 2 vdd
rlabel alu1 541 200 541 200 1 p3
rlabel alu1 562 204 562 204 1 q3
rlabel alu1 554 192 554 192 1 q3
rlabel alu1 534 100 534 100 4 vss
rlabel alu1 534 164 534 164 4 vdd
rlabel alu1 506 152 506 152 1 cnt
rlabel alu1 514 144 514 144 1 cnt
rlabel alu1 562 123 562 123 1 sh0
rlabel alu1 536 132 536 132 1 vss
rlabel alu1 514 120 514 120 1 q1
rlabel alu1 534 92 534 92 2 vss
rlabel alu1 534 28 534 28 2 vdd
rlabel alu1 506 40 506 40 1 cnt
rlabel alu1 514 48 514 48 1 cnt
rlabel alu1 537 59 537 59 1 q0
rlabel alu1 562 67 562 67 1 sh1
rlabel alu1 514 72 514 72 1 q2
rlabel alu1 534 20 534 20 4 vdd
rlabel alu1 534 -44 534 -44 4 vss
rlabel alu1 562 -16 562 -16 1 sh2
rlabel alu1 514 0 514 0 1 cnt
rlabel alu1 506 8 506 8 1 cnt
rlabel alu1 537 -11 537 -11 1 q1
rlabel alu1 514 -24 514 -24 1 q3
rlabel alu1 534 -52 534 -52 2 vss
rlabel alu1 534 -116 534 -116 2 vdd
rlabel alu1 514 -96 514 -96 1 cnt
rlabel alu1 506 -104 506 -104 1 cnt
rlabel alu1 562 -77 562 -77 1 sh3
rlabel alu1 537 -87 537 -87 1 q2
rlabel alu1 516 -72 516 -72 1 vss
<< end >>
